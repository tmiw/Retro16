// from https://github.com/MParygin/v.vga.font8x16
module pc_vga_8x16_00_7F (
		 input		clk,
		 input  [6:0]	ascii_code,
		 input  [3:0]	row,
		 input  [2:0]  col,
		 output wire	row_of_pixels
		 );

reg [255:0] tempval;

always @(posedge clk)
begin
    case (ascii_code[6:1])
		6'h00: tempval <= 256'h00000000000000000000000000000000000000007e818199bd8181a5817e0000;
		6'h01: tempval <= 256'h000000007effffe7c3ffffdbff7e00000000000010387cfefefefe6c00000000;
		6'h02: tempval <= 256'h000000000010387cfe7c381000000000000000003c1818e7e7e73c3c18000000;
		6'h03: tempval <= 256'h000000003c18187effff7e3c18000000000000000000183c3c18000000000000;
		6'h04: tempval <= 256'hffffffffffffe7c3c3e7ffffffffffff00000000003c664242663c0000000000;
		6'h05: tempval <= 256'hffffffffffc399bdbd99c3ffffffffff0000000078cccccccc78321a0e1e0000;
		6'h06: tempval <= 256'h0000000018187e183c666666663c000000000000e0f070303030303f333f0000;
		6'h07: tempval <= 256'h000000c0e6e767636363637f637f0000000000001818db3ce73cdb1818000000;
		6'h08: tempval <= 256'h0000000080c0e0f0f8fef8f0e0c080000000000002060e1e3efe3e1e0e060200;
		6'h09: tempval <= 256'h0000000000183c7e1818187e3c18000000000000666600666666666666660000;
		6'h0A: tempval <= 256'h000000001b1b1b1b1b7bdbdbdb7f00000000007cc60c386cc6c66c3860c67c00;
		6'h0B: tempval <= 256'h00000000fefefefe0000000000000000000000007e183c7e1818187e3c180000;
		6'h0C: tempval <= 256'h00000000181818181818187e3c18000000000000183c7e181818181818180000;
		6'h0D: tempval <= 256'h000000000000180cfe0c1800000000000000000000003060fe60300000000000;
		6'h0E: tempval <= 256'h000000000000fec0c0c00000000000000000000000002466ff66240000000000;
		6'h0F: tempval <= 256'h0000000000fefe7c7c3838100000000000000000001038387c7cfefe00000000;

		6'h10: tempval <= 256'h00000000000000000000000000000000000000001818001818183c3c3c180000;
		6'h11: tempval <= 256'h00000000000000000000002466666600000000006c6cfe6c6c6cfe6c6c000000;
		6'h12: tempval <= 256'h000018187cc68606067cc0c2c67c18180000000086c66030180cc6c200000000;
		6'h13: tempval <= 256'h0000000076ccccccdc76386c6c38000000000000000000000000006030303000;
		6'h14: tempval <= 256'h000000000c18303030303030180c00000000000030180c0c0c0c0c0c18300000;
		6'h15: tempval <= 256'h000000000000663cff3c66000000000000000000000018187e18180000000000;
		6'h16: tempval <= 256'h0000003018181800000000000000000000000000000000007e00000000000000;
		6'h17: tempval <= 256'h000000001818000000000000000000000000000080c06030180c060200000000;
		6'h18: tempval <= 256'h000000007cc6c6e6f6decec6c67c0000000000007e1818181818187838180000;
		6'h19: tempval <= 256'h00000000fec6c06030180c06c67c0000000000007cc60606063c0606c67c0000;
		6'h1A: tempval <= 256'h000000001e0c0c0cfecc6c3c1c0c0000000000007cc6060606fcc0c0c0fe0000;
		6'h1B: tempval <= 256'h000000007cc6c6c6c6fcc0c0603800000000000030303030180c0606c6fe0000;
		6'h1C: tempval <= 256'h000000007cc6c6c6c67cc6c6c67c000000000000780c0606067ec6c6c67c0000;
		6'h1D: tempval <= 256'h0000000000181800000018180000000000000000301818000000181800000000;
		6'h1E: tempval <= 256'h00000000060c18306030180c06000000000000000000007e00007e0000000000;
		6'h1F: tempval <= 256'h000000006030180c060c183060000000000000001818001818180cc6c67c0000;

		6'h20: tempval <= 256'h000000007cc0dcdededec6c6c67c000000000000c6c6c6c6fec6c66c38100000;
		6'h21: tempval <= 256'h00000000fc666666667c666666fc0000000000003c66c2c0c0c0c0c2663c0000;
		6'h22: tempval <= 256'h00000000f86c6666666666666cf8000000000000fe6662606878686266fe0000;
		6'h23: tempval <= 256'h00000000f06060606878686266fe0000000000003a66c6c6dec0c0c2663c0000;
		6'h24: tempval <= 256'h00000000c6c6c6c6c6fec6c6c6c60000000000003c18181818181818183c0000;
		6'h25: tempval <= 256'h0000000078cccccc0c0c0c0c0c1e000000000000e666666c78786c6666e60000;
		6'h26: tempval <= 256'h00000000fe6662606060606060f0000000000000c3c3c3c3c3dbffffe7c30000;
		6'h27: tempval <= 256'h00000000c6c6c6c6cedefef6e6c60000000000007cc6c6c6c6c6c6c6c67c0000;
		6'h28: tempval <= 256'h00000000f0606060607c666666fc000000000e0c7cded6c6c6c6c6c6c67c0000;
		6'h29: tempval <= 256'h00000000e66666666c7c666666fc0000000000007cc6c6060c3860c6c67c0000;
		6'h2A: tempval <= 256'h000000003c18181818181899dbff0000000000007cc6c6c6c6c6c6c6c6c60000;
		6'h2B: tempval <= 256'h00000000183c66c3c3c3c3c3c3c30000000000006666ffdbdbc3c3c3c3c30000;
		6'h2C: tempval <= 256'h00000000c3c3663c18183c66c3c30000000000003c181818183c66c3c3c30000;
		6'h2D: tempval <= 256'h00000000ffc3c16030180c86c3ff0000000000003c30303030303030303c0000;
		6'h2E: tempval <= 256'h0000000002060e1c3870e0c080000000000000003c0c0c0c0c0c0c0c0c3c0000;
		6'h2F: tempval <= 256'h000000000000000000000000c66c38100000ff00000000000000000000000000;
			
			 
		6'h30: tempval <= 256'h000000000000000000000000001830300000000076cccccc7c0c780000000000;
		6'h31: tempval <= 256'h000000007c666666666c786060e00000000000007cc6c0c0c0c67c0000000000;
		6'h32: tempval <= 256'h0000000076cccccccc6c3c0c0c1c0000000000007cc6c0c0fec67c0000000000;
		6'h33: tempval <= 256'h00000000f060606060f060646c3800000078cc0c7ccccccccccc760000000000;
		6'h34: tempval <= 256'h00000000e666666666766c6060e00000000000003c1818181818380018180000;
		6'h35: tempval <= 256'h003c66660606060606060e000606000000000000e6666c78786c666060e00000;
		6'h36: tempval <= 256'h000000003c181818181818181838000000000000dbdbdbdbdbffe60000000000;
		6'h37: tempval <= 256'h00000000666666666666dc0000000000000000007cc6c6c6c6c67c0000000000;
		6'h38: tempval <= 256'h00f060607c6666666666dc0000000000001e0c0c7ccccccccccc760000000000;
		6'h39: tempval <= 256'h00000000f06060606676dc0000000000000000007cc60c3860c67c0000000000;
		6'h3A: tempval <= 256'h000000001c3630303030fc30301000000000000076cccccccccccc0000000000;
		6'h3B: tempval <= 256'h00000000183c66c3c3c3c300000000000000000066ffdbdbc3c3c30000000000;
		6'h3C: tempval <= 256'h00000000c3663c183c66c3000000000000f80c067ec6c6c6c6c6c60000000000;
		6'h3D: tempval <= 256'h00000000fec6603018ccfe0000000000000000000e18181818701818180e0000;
		6'h3E: tempval <= 256'h000000001818181818001818181800000000000070181818180e181818700000;
		6'h3F: tempval <= 256'h000000000000000000000000dc7600000000000000fec6c6c66c381000000000;
	 endcase
end

assign row_of_pixels = tempval[{~ascii_code[0], row, ~col}];
endmodule