// Based on https://github.com/MParygin/v.vga.font8x16
// but converted into a byte-addressed ROM for easier reasoning/management.

module pc_vga_font_rom (
		 input		clk,
		 input  [7:0]	ascii_code,
		 input  [3:0]	row,
		 output reg [7:0]	row_of_pixels
		 );

always @(posedge clk)
begin
    case ({ascii_code, row})
		12'd0: row_of_pixels <= 8'b00000000;
		12'd1: row_of_pixels <= 8'b00000000;
		12'd2: row_of_pixels <= 8'b00000000;
		12'd3: row_of_pixels <= 8'b00000000;
		12'd4: row_of_pixels <= 8'b00000000;
		12'd5: row_of_pixels <= 8'b00000000;
		12'd6: row_of_pixels <= 8'b00000000;
		12'd7: row_of_pixels <= 8'b00000000;
		12'd8: row_of_pixels <= 8'b00000000;
		12'd9: row_of_pixels <= 8'b00000000;
		12'd10: row_of_pixels <= 8'b00000000;
		12'd11: row_of_pixels <= 8'b00000000;
		12'd12: row_of_pixels <= 8'b00000000;
		12'd13: row_of_pixels <= 8'b00000000;
		12'd14: row_of_pixels <= 8'b00000000;
		12'd15: row_of_pixels <= 8'b00000000;
		12'd16: row_of_pixels <= 8'b00000000;
		12'd17: row_of_pixels <= 8'b00000000;
		12'd18: row_of_pixels <= 8'b01111110;
		12'd19: row_of_pixels <= 8'b10000001;
		12'd20: row_of_pixels <= 8'b10100101;
		12'd21: row_of_pixels <= 8'b10000001;
		12'd22: row_of_pixels <= 8'b10000001;
		12'd23: row_of_pixels <= 8'b10111101;
		12'd24: row_of_pixels <= 8'b10011001;
		12'd25: row_of_pixels <= 8'b10000001;
		12'd26: row_of_pixels <= 8'b10000001;
		12'd27: row_of_pixels <= 8'b01111110;
		12'd28: row_of_pixels <= 8'b00000000;
		12'd29: row_of_pixels <= 8'b00000000;
		12'd30: row_of_pixels <= 8'b00000000;
		12'd31: row_of_pixels <= 8'b00000000;
		12'd32: row_of_pixels <= 8'b00000000;
		12'd33: row_of_pixels <= 8'b00000000;
		12'd34: row_of_pixels <= 8'b01111110;
		12'd35: row_of_pixels <= 8'b11111111;
		12'd36: row_of_pixels <= 8'b11011011;
		12'd37: row_of_pixels <= 8'b11111111;
		12'd38: row_of_pixels <= 8'b11111111;
		12'd39: row_of_pixels <= 8'b11000011;
		12'd40: row_of_pixels <= 8'b11100111;
		12'd41: row_of_pixels <= 8'b11111111;
		12'd42: row_of_pixels <= 8'b11111111;
		12'd43: row_of_pixels <= 8'b01111110;
		12'd44: row_of_pixels <= 8'b00000000;
		12'd45: row_of_pixels <= 8'b00000000;
		12'd46: row_of_pixels <= 8'b00000000;
		12'd47: row_of_pixels <= 8'b00000000;
		12'd48: row_of_pixels <= 8'b00000000;
		12'd49: row_of_pixels <= 8'b00000000;
		12'd50: row_of_pixels <= 8'b00000000;
		12'd51: row_of_pixels <= 8'b00000000;
		12'd52: row_of_pixels <= 8'b00110110;
		12'd53: row_of_pixels <= 8'b01111111;
		12'd54: row_of_pixels <= 8'b01111111;
		12'd55: row_of_pixels <= 8'b01111111;
		12'd56: row_of_pixels <= 8'b01111111;
		12'd57: row_of_pixels <= 8'b00111110;
		12'd58: row_of_pixels <= 8'b00011100;
		12'd59: row_of_pixels <= 8'b00001000;
		12'd60: row_of_pixels <= 8'b00000000;
		12'd61: row_of_pixels <= 8'b00000000;
		12'd62: row_of_pixels <= 8'b00000000;
		12'd63: row_of_pixels <= 8'b00000000;
		12'd64: row_of_pixels <= 8'b00000000;
		12'd65: row_of_pixels <= 8'b00000000;
		12'd66: row_of_pixels <= 8'b00000000;
		12'd67: row_of_pixels <= 8'b00000000;
		12'd68: row_of_pixels <= 8'b00001000;
		12'd69: row_of_pixels <= 8'b00011100;
		12'd70: row_of_pixels <= 8'b00111110;
		12'd71: row_of_pixels <= 8'b01111111;
		12'd72: row_of_pixels <= 8'b00111110;
		12'd73: row_of_pixels <= 8'b00011100;
		12'd74: row_of_pixels <= 8'b00001000;
		12'd75: row_of_pixels <= 8'b00000000;
		12'd76: row_of_pixels <= 8'b00000000;
		12'd77: row_of_pixels <= 8'b00000000;
		12'd78: row_of_pixels <= 8'b00000000;
		12'd79: row_of_pixels <= 8'b00000000;
		12'd80: row_of_pixels <= 8'b00000000;
		12'd81: row_of_pixels <= 8'b00000000;
		12'd82: row_of_pixels <= 8'b00000000;
		12'd83: row_of_pixels <= 8'b00011000;
		12'd84: row_of_pixels <= 8'b00111100;
		12'd85: row_of_pixels <= 8'b00111100;
		12'd86: row_of_pixels <= 8'b11100111;
		12'd87: row_of_pixels <= 8'b11100111;
		12'd88: row_of_pixels <= 8'b11100111;
		12'd89: row_of_pixels <= 8'b00011000;
		12'd90: row_of_pixels <= 8'b00011000;
		12'd91: row_of_pixels <= 8'b00111100;
		12'd92: row_of_pixels <= 8'b00000000;
		12'd93: row_of_pixels <= 8'b00000000;
		12'd94: row_of_pixels <= 8'b00000000;
		12'd95: row_of_pixels <= 8'b00000000;
		12'd96: row_of_pixels <= 8'b00000000;
		12'd97: row_of_pixels <= 8'b00000000;
		12'd98: row_of_pixels <= 8'b00000000;
		12'd99: row_of_pixels <= 8'b00011000;
		12'd100: row_of_pixels <= 8'b00111100;
		12'd101: row_of_pixels <= 8'b01111110;
		12'd102: row_of_pixels <= 8'b11111111;
		12'd103: row_of_pixels <= 8'b11111111;
		12'd104: row_of_pixels <= 8'b01111110;
		12'd105: row_of_pixels <= 8'b00011000;
		12'd106: row_of_pixels <= 8'b00011000;
		12'd107: row_of_pixels <= 8'b00111100;
		12'd108: row_of_pixels <= 8'b00000000;
		12'd109: row_of_pixels <= 8'b00000000;
		12'd110: row_of_pixels <= 8'b00000000;
		12'd111: row_of_pixels <= 8'b00000000;
		12'd112: row_of_pixels <= 8'b00000000;
		12'd113: row_of_pixels <= 8'b00000000;
		12'd114: row_of_pixels <= 8'b00000000;
		12'd115: row_of_pixels <= 8'b00000000;
		12'd116: row_of_pixels <= 8'b00000000;
		12'd117: row_of_pixels <= 8'b00000000;
		12'd118: row_of_pixels <= 8'b00011000;
		12'd119: row_of_pixels <= 8'b00111100;
		12'd120: row_of_pixels <= 8'b00111100;
		12'd121: row_of_pixels <= 8'b00011000;
		12'd122: row_of_pixels <= 8'b00000000;
		12'd123: row_of_pixels <= 8'b00000000;
		12'd124: row_of_pixels <= 8'b00000000;
		12'd125: row_of_pixels <= 8'b00000000;
		12'd126: row_of_pixels <= 8'b00000000;
		12'd127: row_of_pixels <= 8'b00000000;
		12'd128: row_of_pixels <= 8'b11111111;
		12'd129: row_of_pixels <= 8'b11111111;
		12'd130: row_of_pixels <= 8'b11111111;
		12'd131: row_of_pixels <= 8'b11111111;
		12'd132: row_of_pixels <= 8'b11111111;
		12'd133: row_of_pixels <= 8'b11111111;
		12'd134: row_of_pixels <= 8'b11100111;
		12'd135: row_of_pixels <= 8'b11000011;
		12'd136: row_of_pixels <= 8'b11000011;
		12'd137: row_of_pixels <= 8'b11100111;
		12'd138: row_of_pixels <= 8'b11111111;
		12'd139: row_of_pixels <= 8'b11111111;
		12'd140: row_of_pixels <= 8'b11111111;
		12'd141: row_of_pixels <= 8'b11111111;
		12'd142: row_of_pixels <= 8'b11111111;
		12'd143: row_of_pixels <= 8'b11111111;
		12'd144: row_of_pixels <= 8'b00000000;
		12'd145: row_of_pixels <= 8'b00000000;
		12'd146: row_of_pixels <= 8'b00000000;
		12'd147: row_of_pixels <= 8'b00000000;
		12'd148: row_of_pixels <= 8'b00000000;
		12'd149: row_of_pixels <= 8'b00111100;
		12'd150: row_of_pixels <= 8'b01100110;
		12'd151: row_of_pixels <= 8'b01000010;
		12'd152: row_of_pixels <= 8'b01000010;
		12'd153: row_of_pixels <= 8'b01100110;
		12'd154: row_of_pixels <= 8'b00111100;
		12'd155: row_of_pixels <= 8'b00000000;
		12'd156: row_of_pixels <= 8'b00000000;
		12'd157: row_of_pixels <= 8'b00000000;
		12'd158: row_of_pixels <= 8'b00000000;
		12'd159: row_of_pixels <= 8'b00000000;
		12'd160: row_of_pixels <= 8'b11111111;
		12'd161: row_of_pixels <= 8'b11111111;
		12'd162: row_of_pixels <= 8'b11111111;
		12'd163: row_of_pixels <= 8'b11111111;
		12'd164: row_of_pixels <= 8'b11111111;
		12'd165: row_of_pixels <= 8'b11000011;
		12'd166: row_of_pixels <= 8'b10011001;
		12'd167: row_of_pixels <= 8'b10111101;
		12'd168: row_of_pixels <= 8'b10111101;
		12'd169: row_of_pixels <= 8'b10011001;
		12'd170: row_of_pixels <= 8'b11000011;
		12'd171: row_of_pixels <= 8'b11111111;
		12'd172: row_of_pixels <= 8'b11111111;
		12'd173: row_of_pixels <= 8'b11111111;
		12'd174: row_of_pixels <= 8'b11111111;
		12'd175: row_of_pixels <= 8'b11111111;
		12'd176: row_of_pixels <= 8'b00000000;
		12'd177: row_of_pixels <= 8'b00000000;
		12'd178: row_of_pixels <= 8'b01111000;
		12'd179: row_of_pixels <= 8'b01110000;
		12'd180: row_of_pixels <= 8'b01011000;
		12'd181: row_of_pixels <= 8'b01001100;
		12'd182: row_of_pixels <= 8'b00011110;
		12'd183: row_of_pixels <= 8'b00110011;
		12'd184: row_of_pixels <= 8'b00110011;
		12'd185: row_of_pixels <= 8'b00110011;
		12'd186: row_of_pixels <= 8'b00110011;
		12'd187: row_of_pixels <= 8'b00011110;
		12'd188: row_of_pixels <= 8'b00000000;
		12'd189: row_of_pixels <= 8'b00000000;
		12'd190: row_of_pixels <= 8'b00000000;
		12'd191: row_of_pixels <= 8'b00000000;
		12'd192: row_of_pixels <= 8'b00000000;
		12'd193: row_of_pixels <= 8'b00000000;
		12'd194: row_of_pixels <= 8'b00111100;
		12'd195: row_of_pixels <= 8'b01100110;
		12'd196: row_of_pixels <= 8'b01100110;
		12'd197: row_of_pixels <= 8'b01100110;
		12'd198: row_of_pixels <= 8'b01100110;
		12'd199: row_of_pixels <= 8'b00111100;
		12'd200: row_of_pixels <= 8'b00011000;
		12'd201: row_of_pixels <= 8'b01111110;
		12'd202: row_of_pixels <= 8'b00011000;
		12'd203: row_of_pixels <= 8'b00011000;
		12'd204: row_of_pixels <= 8'b00000000;
		12'd205: row_of_pixels <= 8'b00000000;
		12'd206: row_of_pixels <= 8'b00000000;
		12'd207: row_of_pixels <= 8'b00000000;
		12'd208: row_of_pixels <= 8'b00000000;
		12'd209: row_of_pixels <= 8'b00000000;
		12'd210: row_of_pixels <= 8'b11111100;
		12'd211: row_of_pixels <= 8'b11001100;
		12'd212: row_of_pixels <= 8'b11111100;
		12'd213: row_of_pixels <= 8'b00001100;
		12'd214: row_of_pixels <= 8'b00001100;
		12'd215: row_of_pixels <= 8'b00001100;
		12'd216: row_of_pixels <= 8'b00001100;
		12'd217: row_of_pixels <= 8'b00001110;
		12'd218: row_of_pixels <= 8'b00001111;
		12'd219: row_of_pixels <= 8'b00000111;
		12'd220: row_of_pixels <= 8'b00000000;
		12'd221: row_of_pixels <= 8'b00000000;
		12'd222: row_of_pixels <= 8'b00000000;
		12'd223: row_of_pixels <= 8'b00000000;
		12'd224: row_of_pixels <= 8'b00000000;
		12'd225: row_of_pixels <= 8'b00000000;
		12'd226: row_of_pixels <= 8'b11111110;
		12'd227: row_of_pixels <= 8'b11000110;
		12'd228: row_of_pixels <= 8'b11111110;
		12'd229: row_of_pixels <= 8'b11000110;
		12'd230: row_of_pixels <= 8'b11000110;
		12'd231: row_of_pixels <= 8'b11000110;
		12'd232: row_of_pixels <= 8'b11000110;
		12'd233: row_of_pixels <= 8'b11100110;
		12'd234: row_of_pixels <= 8'b11100111;
		12'd235: row_of_pixels <= 8'b01100111;
		12'd236: row_of_pixels <= 8'b00000011;
		12'd237: row_of_pixels <= 8'b00000000;
		12'd238: row_of_pixels <= 8'b00000000;
		12'd239: row_of_pixels <= 8'b00000000;
		12'd240: row_of_pixels <= 8'b00000000;
		12'd241: row_of_pixels <= 8'b00000000;
		12'd242: row_of_pixels <= 8'b00000000;
		12'd243: row_of_pixels <= 8'b00011000;
		12'd244: row_of_pixels <= 8'b00011000;
		12'd245: row_of_pixels <= 8'b11011011;
		12'd246: row_of_pixels <= 8'b00111100;
		12'd247: row_of_pixels <= 8'b11100111;
		12'd248: row_of_pixels <= 8'b00111100;
		12'd249: row_of_pixels <= 8'b11011011;
		12'd250: row_of_pixels <= 8'b00011000;
		12'd251: row_of_pixels <= 8'b00011000;
		12'd252: row_of_pixels <= 8'b00000000;
		12'd253: row_of_pixels <= 8'b00000000;
		12'd254: row_of_pixels <= 8'b00000000;
		12'd255: row_of_pixels <= 8'b00000000;
		12'd256: row_of_pixels <= 8'b00000000;
		12'd257: row_of_pixels <= 8'b00000001;
		12'd258: row_of_pixels <= 8'b00000011;
		12'd259: row_of_pixels <= 8'b00000111;
		12'd260: row_of_pixels <= 8'b00001111;
		12'd261: row_of_pixels <= 8'b00011111;
		12'd262: row_of_pixels <= 8'b01111111;
		12'd263: row_of_pixels <= 8'b00011111;
		12'd264: row_of_pixels <= 8'b00001111;
		12'd265: row_of_pixels <= 8'b00000111;
		12'd266: row_of_pixels <= 8'b00000011;
		12'd267: row_of_pixels <= 8'b00000001;
		12'd268: row_of_pixels <= 8'b00000000;
		12'd269: row_of_pixels <= 8'b00000000;
		12'd270: row_of_pixels <= 8'b00000000;
		12'd271: row_of_pixels <= 8'b00000000;
		12'd272: row_of_pixels <= 8'b00000000;
		12'd273: row_of_pixels <= 8'b01000000;
		12'd274: row_of_pixels <= 8'b01100000;
		12'd275: row_of_pixels <= 8'b01110000;
		12'd276: row_of_pixels <= 8'b01111000;
		12'd277: row_of_pixels <= 8'b01111100;
		12'd278: row_of_pixels <= 8'b01111111;
		12'd279: row_of_pixels <= 8'b01111100;
		12'd280: row_of_pixels <= 8'b01111000;
		12'd281: row_of_pixels <= 8'b01110000;
		12'd282: row_of_pixels <= 8'b01100000;
		12'd283: row_of_pixels <= 8'b01000000;
		12'd284: row_of_pixels <= 8'b00000000;
		12'd285: row_of_pixels <= 8'b00000000;
		12'd286: row_of_pixels <= 8'b00000000;
		12'd287: row_of_pixels <= 8'b00000000;
		12'd288: row_of_pixels <= 8'b00000000;
		12'd289: row_of_pixels <= 8'b00000000;
		12'd290: row_of_pixels <= 8'b00011000;
		12'd291: row_of_pixels <= 8'b00111100;
		12'd292: row_of_pixels <= 8'b01111110;
		12'd293: row_of_pixels <= 8'b00011000;
		12'd294: row_of_pixels <= 8'b00011000;
		12'd295: row_of_pixels <= 8'b00011000;
		12'd296: row_of_pixels <= 8'b01111110;
		12'd297: row_of_pixels <= 8'b00111100;
		12'd298: row_of_pixels <= 8'b00011000;
		12'd299: row_of_pixels <= 8'b00000000;
		12'd300: row_of_pixels <= 8'b00000000;
		12'd301: row_of_pixels <= 8'b00000000;
		12'd302: row_of_pixels <= 8'b00000000;
		12'd303: row_of_pixels <= 8'b00000000;
		12'd304: row_of_pixels <= 8'b00000000;
		12'd305: row_of_pixels <= 8'b00000000;
		12'd306: row_of_pixels <= 8'b01100110;
		12'd307: row_of_pixels <= 8'b01100110;
		12'd308: row_of_pixels <= 8'b01100110;
		12'd309: row_of_pixels <= 8'b01100110;
		12'd310: row_of_pixels <= 8'b01100110;
		12'd311: row_of_pixels <= 8'b01100110;
		12'd312: row_of_pixels <= 8'b01100110;
		12'd313: row_of_pixels <= 8'b00000000;
		12'd314: row_of_pixels <= 8'b01100110;
		12'd315: row_of_pixels <= 8'b01100110;
		12'd316: row_of_pixels <= 8'b00000000;
		12'd317: row_of_pixels <= 8'b00000000;
		12'd318: row_of_pixels <= 8'b00000000;
		12'd319: row_of_pixels <= 8'b00000000;
		12'd320: row_of_pixels <= 8'b00000000;
		12'd321: row_of_pixels <= 8'b00000000;
		12'd322: row_of_pixels <= 8'b11111110;
		12'd323: row_of_pixels <= 8'b11011011;
		12'd324: row_of_pixels <= 8'b11011011;
		12'd325: row_of_pixels <= 8'b11011011;
		12'd326: row_of_pixels <= 8'b11011110;
		12'd327: row_of_pixels <= 8'b11011000;
		12'd328: row_of_pixels <= 8'b11011000;
		12'd329: row_of_pixels <= 8'b11011000;
		12'd330: row_of_pixels <= 8'b11011000;
		12'd331: row_of_pixels <= 8'b11011000;
		12'd332: row_of_pixels <= 8'b00000000;
		12'd333: row_of_pixels <= 8'b00000000;
		12'd334: row_of_pixels <= 8'b00000000;
		12'd335: row_of_pixels <= 8'b00000000;
		12'd336: row_of_pixels <= 8'b00000000;
		12'd337: row_of_pixels <= 8'b00111110;
		12'd338: row_of_pixels <= 8'b01100011;
		12'd339: row_of_pixels <= 8'b00000110;
		12'd340: row_of_pixels <= 8'b00011100;
		12'd341: row_of_pixels <= 8'b00110110;
		12'd342: row_of_pixels <= 8'b01100011;
		12'd343: row_of_pixels <= 8'b01100011;
		12'd344: row_of_pixels <= 8'b00110110;
		12'd345: row_of_pixels <= 8'b00011100;
		12'd346: row_of_pixels <= 8'b00110000;
		12'd347: row_of_pixels <= 8'b01100011;
		12'd348: row_of_pixels <= 8'b00111110;
		12'd349: row_of_pixels <= 8'b00000000;
		12'd350: row_of_pixels <= 8'b00000000;
		12'd351: row_of_pixels <= 8'b00000000;
		12'd352: row_of_pixels <= 8'b00000000;
		12'd353: row_of_pixels <= 8'b00000000;
		12'd354: row_of_pixels <= 8'b00000000;
		12'd355: row_of_pixels <= 8'b00000000;
		12'd356: row_of_pixels <= 8'b00000000;
		12'd357: row_of_pixels <= 8'b00000000;
		12'd358: row_of_pixels <= 8'b00000000;
		12'd359: row_of_pixels <= 8'b00000000;
		12'd360: row_of_pixels <= 8'b01111111;
		12'd361: row_of_pixels <= 8'b01111111;
		12'd362: row_of_pixels <= 8'b01111111;
		12'd363: row_of_pixels <= 8'b01111111;
		12'd364: row_of_pixels <= 8'b00000000;
		12'd365: row_of_pixels <= 8'b00000000;
		12'd366: row_of_pixels <= 8'b00000000;
		12'd367: row_of_pixels <= 8'b00000000;
		12'd368: row_of_pixels <= 8'b00000000;
		12'd369: row_of_pixels <= 8'b00000000;
		12'd370: row_of_pixels <= 8'b00011000;
		12'd371: row_of_pixels <= 8'b00111100;
		12'd372: row_of_pixels <= 8'b01111110;
		12'd373: row_of_pixels <= 8'b00011000;
		12'd374: row_of_pixels <= 8'b00011000;
		12'd375: row_of_pixels <= 8'b00011000;
		12'd376: row_of_pixels <= 8'b01111110;
		12'd377: row_of_pixels <= 8'b00111100;
		12'd378: row_of_pixels <= 8'b00011000;
		12'd379: row_of_pixels <= 8'b01111110;
		12'd380: row_of_pixels <= 8'b00000000;
		12'd381: row_of_pixels <= 8'b00000000;
		12'd382: row_of_pixels <= 8'b00000000;
		12'd383: row_of_pixels <= 8'b00000000;
		12'd384: row_of_pixels <= 8'b00000000;
		12'd385: row_of_pixels <= 8'b00000000;
		12'd386: row_of_pixels <= 8'b00011000;
		12'd387: row_of_pixels <= 8'b00111100;
		12'd388: row_of_pixels <= 8'b01111110;
		12'd389: row_of_pixels <= 8'b00011000;
		12'd390: row_of_pixels <= 8'b00011000;
		12'd391: row_of_pixels <= 8'b00011000;
		12'd392: row_of_pixels <= 8'b00011000;
		12'd393: row_of_pixels <= 8'b00011000;
		12'd394: row_of_pixels <= 8'b00011000;
		12'd395: row_of_pixels <= 8'b00011000;
		12'd396: row_of_pixels <= 8'b00000000;
		12'd397: row_of_pixels <= 8'b00000000;
		12'd398: row_of_pixels <= 8'b00000000;
		12'd399: row_of_pixels <= 8'b00000000;
		12'd400: row_of_pixels <= 8'b00000000;
		12'd401: row_of_pixels <= 8'b00000000;
		12'd402: row_of_pixels <= 8'b00011000;
		12'd403: row_of_pixels <= 8'b00011000;
		12'd404: row_of_pixels <= 8'b00011000;
		12'd405: row_of_pixels <= 8'b00011000;
		12'd406: row_of_pixels <= 8'b00011000;
		12'd407: row_of_pixels <= 8'b00011000;
		12'd408: row_of_pixels <= 8'b00011000;
		12'd409: row_of_pixels <= 8'b01111110;
		12'd410: row_of_pixels <= 8'b00111100;
		12'd411: row_of_pixels <= 8'b00011000;
		12'd412: row_of_pixels <= 8'b00000000;
		12'd413: row_of_pixels <= 8'b00000000;
		12'd414: row_of_pixels <= 8'b00000000;
		12'd415: row_of_pixels <= 8'b00000000;
		12'd416: row_of_pixels <= 8'b00000000;
		12'd417: row_of_pixels <= 8'b00000000;
		12'd418: row_of_pixels <= 8'b00000000;
		12'd419: row_of_pixels <= 8'b00000000;
		12'd420: row_of_pixels <= 8'b00000000;
		12'd421: row_of_pixels <= 8'b00011000;
		12'd422: row_of_pixels <= 8'b00110000;
		12'd423: row_of_pixels <= 8'b01111111;
		12'd424: row_of_pixels <= 8'b00110000;
		12'd425: row_of_pixels <= 8'b00011000;
		12'd426: row_of_pixels <= 8'b00000000;
		12'd427: row_of_pixels <= 8'b00000000;
		12'd428: row_of_pixels <= 8'b00000000;
		12'd429: row_of_pixels <= 8'b00000000;
		12'd430: row_of_pixels <= 8'b00000000;
		12'd431: row_of_pixels <= 8'b00000000;
		12'd432: row_of_pixels <= 8'b00000000;
		12'd433: row_of_pixels <= 8'b00000000;
		12'd434: row_of_pixels <= 8'b00000000;
		12'd435: row_of_pixels <= 8'b00000000;
		12'd436: row_of_pixels <= 8'b00000000;
		12'd437: row_of_pixels <= 8'b00001100;
		12'd438: row_of_pixels <= 8'b00000110;
		12'd439: row_of_pixels <= 8'b01111111;
		12'd440: row_of_pixels <= 8'b00000110;
		12'd441: row_of_pixels <= 8'b00001100;
		12'd442: row_of_pixels <= 8'b00000000;
		12'd443: row_of_pixels <= 8'b00000000;
		12'd444: row_of_pixels <= 8'b00000000;
		12'd445: row_of_pixels <= 8'b00000000;
		12'd446: row_of_pixels <= 8'b00000000;
		12'd447: row_of_pixels <= 8'b00000000;
		12'd448: row_of_pixels <= 8'b00000000;
		12'd449: row_of_pixels <= 8'b00000000;
		12'd450: row_of_pixels <= 8'b00000000;
		12'd451: row_of_pixels <= 8'b00000000;
		12'd452: row_of_pixels <= 8'b00000000;
		12'd453: row_of_pixels <= 8'b00000000;
		12'd454: row_of_pixels <= 8'b00000011;
		12'd455: row_of_pixels <= 8'b00000011;
		12'd456: row_of_pixels <= 8'b00000011;
		12'd457: row_of_pixels <= 8'b01111111;
		12'd458: row_of_pixels <= 8'b00000000;
		12'd459: row_of_pixels <= 8'b00000000;
		12'd460: row_of_pixels <= 8'b00000000;
		12'd461: row_of_pixels <= 8'b00000000;
		12'd462: row_of_pixels <= 8'b00000000;
		12'd463: row_of_pixels <= 8'b00000000;
		12'd464: row_of_pixels <= 8'b00000000;
		12'd465: row_of_pixels <= 8'b00000000;
		12'd466: row_of_pixels <= 8'b00000000;
		12'd467: row_of_pixels <= 8'b00000000;
		12'd468: row_of_pixels <= 8'b00000000;
		12'd469: row_of_pixels <= 8'b00100100;
		12'd470: row_of_pixels <= 8'b01100110;
		12'd471: row_of_pixels <= 8'b11111111;
		12'd472: row_of_pixels <= 8'b01100110;
		12'd473: row_of_pixels <= 8'b00100100;
		12'd474: row_of_pixels <= 8'b00000000;
		12'd475: row_of_pixels <= 8'b00000000;
		12'd476: row_of_pixels <= 8'b00000000;
		12'd477: row_of_pixels <= 8'b00000000;
		12'd478: row_of_pixels <= 8'b00000000;
		12'd479: row_of_pixels <= 8'b00000000;
		12'd480: row_of_pixels <= 8'b00000000;
		12'd481: row_of_pixels <= 8'b00000000;
		12'd482: row_of_pixels <= 8'b00000000;
		12'd483: row_of_pixels <= 8'b00000000;
		12'd484: row_of_pixels <= 8'b00001000;
		12'd485: row_of_pixels <= 8'b00011100;
		12'd486: row_of_pixels <= 8'b00011100;
		12'd487: row_of_pixels <= 8'b00111110;
		12'd488: row_of_pixels <= 8'b00111110;
		12'd489: row_of_pixels <= 8'b01111111;
		12'd490: row_of_pixels <= 8'b01111111;
		12'd491: row_of_pixels <= 8'b00000000;
		12'd492: row_of_pixels <= 8'b00000000;
		12'd493: row_of_pixels <= 8'b00000000;
		12'd494: row_of_pixels <= 8'b00000000;
		12'd495: row_of_pixels <= 8'b00000000;
		12'd496: row_of_pixels <= 8'b00000000;
		12'd497: row_of_pixels <= 8'b00000000;
		12'd498: row_of_pixels <= 8'b00000000;
		12'd499: row_of_pixels <= 8'b00000000;
		12'd500: row_of_pixels <= 8'b01111111;
		12'd501: row_of_pixels <= 8'b01111111;
		12'd502: row_of_pixels <= 8'b00111110;
		12'd503: row_of_pixels <= 8'b00111110;
		12'd504: row_of_pixels <= 8'b00011100;
		12'd505: row_of_pixels <= 8'b00011100;
		12'd506: row_of_pixels <= 8'b00001000;
		12'd507: row_of_pixels <= 8'b00000000;
		12'd508: row_of_pixels <= 8'b00000000;
		12'd509: row_of_pixels <= 8'b00000000;
		12'd510: row_of_pixels <= 8'b00000000;
		12'd511: row_of_pixels <= 8'b00000000;
		12'd512: row_of_pixels <= 8'b00000000;
		12'd513: row_of_pixels <= 8'b00000000;
		12'd514: row_of_pixels <= 8'b00000000;
		12'd515: row_of_pixels <= 8'b00000000;
		12'd516: row_of_pixels <= 8'b00000000;
		12'd517: row_of_pixels <= 8'b00000000;
		12'd518: row_of_pixels <= 8'b00000000;
		12'd519: row_of_pixels <= 8'b00000000;
		12'd520: row_of_pixels <= 8'b00000000;
		12'd521: row_of_pixels <= 8'b00000000;
		12'd522: row_of_pixels <= 8'b00000000;
		12'd523: row_of_pixels <= 8'b00000000;
		12'd524: row_of_pixels <= 8'b00000000;
		12'd525: row_of_pixels <= 8'b00000000;
		12'd526: row_of_pixels <= 8'b00000000;
		12'd527: row_of_pixels <= 8'b00000000;
		12'd528: row_of_pixels <= 8'b00000000;
		12'd529: row_of_pixels <= 8'b00000000;
		12'd530: row_of_pixels <= 8'b00011000;
		12'd531: row_of_pixels <= 8'b00111100;
		12'd532: row_of_pixels <= 8'b00111100;
		12'd533: row_of_pixels <= 8'b00111100;
		12'd534: row_of_pixels <= 8'b00011000;
		12'd535: row_of_pixels <= 8'b00011000;
		12'd536: row_of_pixels <= 8'b00011000;
		12'd537: row_of_pixels <= 8'b00000000;
		12'd538: row_of_pixels <= 8'b00011000;
		12'd539: row_of_pixels <= 8'b00011000;
		12'd540: row_of_pixels <= 8'b00000000;
		12'd541: row_of_pixels <= 8'b00000000;
		12'd542: row_of_pixels <= 8'b00000000;
		12'd543: row_of_pixels <= 8'b00000000;
		12'd544: row_of_pixels <= 8'b00000000;
		12'd545: row_of_pixels <= 8'b01100110;
		12'd546: row_of_pixels <= 8'b01100110;
		12'd547: row_of_pixels <= 8'b01100110;
		12'd548: row_of_pixels <= 8'b00100100;
		12'd549: row_of_pixels <= 8'b00000000;
		12'd550: row_of_pixels <= 8'b00000000;
		12'd551: row_of_pixels <= 8'b00000000;
		12'd552: row_of_pixels <= 8'b00000000;
		12'd553: row_of_pixels <= 8'b00000000;
		12'd554: row_of_pixels <= 8'b00000000;
		12'd555: row_of_pixels <= 8'b00000000;
		12'd556: row_of_pixels <= 8'b00000000;
		12'd557: row_of_pixels <= 8'b00000000;
		12'd558: row_of_pixels <= 8'b00000000;
		12'd559: row_of_pixels <= 8'b00000000;
		12'd560: row_of_pixels <= 8'b00000000;
		12'd561: row_of_pixels <= 8'b00000000;
		12'd562: row_of_pixels <= 8'b00000000;
		12'd563: row_of_pixels <= 8'b00110110;
		12'd564: row_of_pixels <= 8'b00110110;
		12'd565: row_of_pixels <= 8'b01111111;
		12'd566: row_of_pixels <= 8'b00110110;
		12'd567: row_of_pixels <= 8'b00110110;
		12'd568: row_of_pixels <= 8'b00110110;
		12'd569: row_of_pixels <= 8'b01111111;
		12'd570: row_of_pixels <= 8'b00110110;
		12'd571: row_of_pixels <= 8'b00110110;
		12'd572: row_of_pixels <= 8'b00000000;
		12'd573: row_of_pixels <= 8'b00000000;
		12'd574: row_of_pixels <= 8'b00000000;
		12'd575: row_of_pixels <= 8'b00000000;
		12'd576: row_of_pixels <= 8'b00011000;
		12'd577: row_of_pixels <= 8'b00011000;
		12'd578: row_of_pixels <= 8'b00111110;
		12'd579: row_of_pixels <= 8'b01100011;
		12'd580: row_of_pixels <= 8'b01000011;
		12'd581: row_of_pixels <= 8'b00000011;
		12'd582: row_of_pixels <= 8'b00111110;
		12'd583: row_of_pixels <= 8'b01100000;
		12'd584: row_of_pixels <= 8'b01100000;
		12'd585: row_of_pixels <= 8'b01100001;
		12'd586: row_of_pixels <= 8'b01100011;
		12'd587: row_of_pixels <= 8'b00111110;
		12'd588: row_of_pixels <= 8'b00011000;
		12'd589: row_of_pixels <= 8'b00011000;
		12'd590: row_of_pixels <= 8'b00000000;
		12'd591: row_of_pixels <= 8'b00000000;
		12'd592: row_of_pixels <= 8'b00000000;
		12'd593: row_of_pixels <= 8'b00000000;
		12'd594: row_of_pixels <= 8'b00000000;
		12'd595: row_of_pixels <= 8'b00000000;
		12'd596: row_of_pixels <= 8'b01000011;
		12'd597: row_of_pixels <= 8'b01100011;
		12'd598: row_of_pixels <= 8'b00110000;
		12'd599: row_of_pixels <= 8'b00011000;
		12'd600: row_of_pixels <= 8'b00001100;
		12'd601: row_of_pixels <= 8'b00000110;
		12'd602: row_of_pixels <= 8'b01100011;
		12'd603: row_of_pixels <= 8'b01100001;
		12'd604: row_of_pixels <= 8'b00000000;
		12'd605: row_of_pixels <= 8'b00000000;
		12'd606: row_of_pixels <= 8'b00000000;
		12'd607: row_of_pixels <= 8'b00000000;
		12'd608: row_of_pixels <= 8'b00000000;
		12'd609: row_of_pixels <= 8'b00000000;
		12'd610: row_of_pixels <= 8'b00011100;
		12'd611: row_of_pixels <= 8'b00110110;
		12'd612: row_of_pixels <= 8'b00110110;
		12'd613: row_of_pixels <= 8'b00011100;
		12'd614: row_of_pixels <= 8'b01101110;
		12'd615: row_of_pixels <= 8'b00111011;
		12'd616: row_of_pixels <= 8'b00110011;
		12'd617: row_of_pixels <= 8'b00110011;
		12'd618: row_of_pixels <= 8'b00110011;
		12'd619: row_of_pixels <= 8'b01101110;
		12'd620: row_of_pixels <= 8'b00000000;
		12'd621: row_of_pixels <= 8'b00000000;
		12'd622: row_of_pixels <= 8'b00000000;
		12'd623: row_of_pixels <= 8'b00000000;
		12'd624: row_of_pixels <= 8'b00000000;
		12'd625: row_of_pixels <= 8'b00001100;
		12'd626: row_of_pixels <= 8'b00001100;
		12'd627: row_of_pixels <= 8'b00001100;
		12'd628: row_of_pixels <= 8'b00000110;
		12'd629: row_of_pixels <= 8'b00000000;
		12'd630: row_of_pixels <= 8'b00000000;
		12'd631: row_of_pixels <= 8'b00000000;
		12'd632: row_of_pixels <= 8'b00000000;
		12'd633: row_of_pixels <= 8'b00000000;
		12'd634: row_of_pixels <= 8'b00000000;
		12'd635: row_of_pixels <= 8'b00000000;
		12'd636: row_of_pixels <= 8'b00000000;
		12'd637: row_of_pixels <= 8'b00000000;
		12'd638: row_of_pixels <= 8'b00000000;
		12'd639: row_of_pixels <= 8'b00000000;
		12'd640: row_of_pixels <= 8'b00000000;
		12'd641: row_of_pixels <= 8'b00000000;
		12'd642: row_of_pixels <= 8'b00110000;
		12'd643: row_of_pixels <= 8'b00011000;
		12'd644: row_of_pixels <= 8'b00001100;
		12'd645: row_of_pixels <= 8'b00001100;
		12'd646: row_of_pixels <= 8'b00001100;
		12'd647: row_of_pixels <= 8'b00001100;
		12'd648: row_of_pixels <= 8'b00001100;
		12'd649: row_of_pixels <= 8'b00001100;
		12'd650: row_of_pixels <= 8'b00011000;
		12'd651: row_of_pixels <= 8'b00110000;
		12'd652: row_of_pixels <= 8'b00000000;
		12'd653: row_of_pixels <= 8'b00000000;
		12'd654: row_of_pixels <= 8'b00000000;
		12'd655: row_of_pixels <= 8'b00000000;
		12'd656: row_of_pixels <= 8'b00000000;
		12'd657: row_of_pixels <= 8'b00000000;
		12'd658: row_of_pixels <= 8'b00001100;
		12'd659: row_of_pixels <= 8'b00011000;
		12'd660: row_of_pixels <= 8'b00110000;
		12'd661: row_of_pixels <= 8'b00110000;
		12'd662: row_of_pixels <= 8'b00110000;
		12'd663: row_of_pixels <= 8'b00110000;
		12'd664: row_of_pixels <= 8'b00110000;
		12'd665: row_of_pixels <= 8'b00110000;
		12'd666: row_of_pixels <= 8'b00011000;
		12'd667: row_of_pixels <= 8'b00001100;
		12'd668: row_of_pixels <= 8'b00000000;
		12'd669: row_of_pixels <= 8'b00000000;
		12'd670: row_of_pixels <= 8'b00000000;
		12'd671: row_of_pixels <= 8'b00000000;
		12'd672: row_of_pixels <= 8'b00000000;
		12'd673: row_of_pixels <= 8'b00000000;
		12'd674: row_of_pixels <= 8'b00000000;
		12'd675: row_of_pixels <= 8'b00000000;
		12'd676: row_of_pixels <= 8'b00000000;
		12'd677: row_of_pixels <= 8'b01100110;
		12'd678: row_of_pixels <= 8'b00111100;
		12'd679: row_of_pixels <= 8'b11111111;
		12'd680: row_of_pixels <= 8'b00111100;
		12'd681: row_of_pixels <= 8'b01100110;
		12'd682: row_of_pixels <= 8'b00000000;
		12'd683: row_of_pixels <= 8'b00000000;
		12'd684: row_of_pixels <= 8'b00000000;
		12'd685: row_of_pixels <= 8'b00000000;
		12'd686: row_of_pixels <= 8'b00000000;
		12'd687: row_of_pixels <= 8'b00000000;
		12'd688: row_of_pixels <= 8'b00000000;
		12'd689: row_of_pixels <= 8'b00000000;
		12'd690: row_of_pixels <= 8'b00000000;
		12'd691: row_of_pixels <= 8'b00000000;
		12'd692: row_of_pixels <= 8'b00000000;
		12'd693: row_of_pixels <= 8'b00011000;
		12'd694: row_of_pixels <= 8'b00011000;
		12'd695: row_of_pixels <= 8'b01111110;
		12'd696: row_of_pixels <= 8'b00011000;
		12'd697: row_of_pixels <= 8'b00011000;
		12'd698: row_of_pixels <= 8'b00000000;
		12'd699: row_of_pixels <= 8'b00000000;
		12'd700: row_of_pixels <= 8'b00000000;
		12'd701: row_of_pixels <= 8'b00000000;
		12'd702: row_of_pixels <= 8'b00000000;
		12'd703: row_of_pixels <= 8'b00000000;
		12'd704: row_of_pixels <= 8'b00000000;
		12'd705: row_of_pixels <= 8'b00000000;
		12'd706: row_of_pixels <= 8'b00000000;
		12'd707: row_of_pixels <= 8'b00000000;
		12'd708: row_of_pixels <= 8'b00000000;
		12'd709: row_of_pixels <= 8'b00000000;
		12'd710: row_of_pixels <= 8'b00000000;
		12'd711: row_of_pixels <= 8'b00000000;
		12'd712: row_of_pixels <= 8'b00000000;
		12'd713: row_of_pixels <= 8'b00011000;
		12'd714: row_of_pixels <= 8'b00011000;
		12'd715: row_of_pixels <= 8'b00011000;
		12'd716: row_of_pixels <= 8'b00001100;
		12'd717: row_of_pixels <= 8'b00000000;
		12'd718: row_of_pixels <= 8'b00000000;
		12'd719: row_of_pixels <= 8'b00000000;
		12'd720: row_of_pixels <= 8'b00000000;
		12'd721: row_of_pixels <= 8'b00000000;
		12'd722: row_of_pixels <= 8'b00000000;
		12'd723: row_of_pixels <= 8'b00000000;
		12'd724: row_of_pixels <= 8'b00000000;
		12'd725: row_of_pixels <= 8'b00000000;
		12'd726: row_of_pixels <= 8'b00000000;
		12'd727: row_of_pixels <= 8'b01111110;
		12'd728: row_of_pixels <= 8'b00000000;
		12'd729: row_of_pixels <= 8'b00000000;
		12'd730: row_of_pixels <= 8'b00000000;
		12'd731: row_of_pixels <= 8'b00000000;
		12'd732: row_of_pixels <= 8'b00000000;
		12'd733: row_of_pixels <= 8'b00000000;
		12'd734: row_of_pixels <= 8'b00000000;
		12'd735: row_of_pixels <= 8'b00000000;
		12'd736: row_of_pixels <= 8'b00000000;
		12'd737: row_of_pixels <= 8'b00000000;
		12'd738: row_of_pixels <= 8'b00000000;
		12'd739: row_of_pixels <= 8'b00000000;
		12'd740: row_of_pixels <= 8'b00000000;
		12'd741: row_of_pixels <= 8'b00000000;
		12'd742: row_of_pixels <= 8'b00000000;
		12'd743: row_of_pixels <= 8'b00000000;
		12'd744: row_of_pixels <= 8'b00000000;
		12'd745: row_of_pixels <= 8'b00000000;
		12'd746: row_of_pixels <= 8'b00011000;
		12'd747: row_of_pixels <= 8'b00011000;
		12'd748: row_of_pixels <= 8'b00000000;
		12'd749: row_of_pixels <= 8'b00000000;
		12'd750: row_of_pixels <= 8'b00000000;
		12'd751: row_of_pixels <= 8'b00000000;
		12'd752: row_of_pixels <= 8'b00000000;
		12'd753: row_of_pixels <= 8'b00000000;
		12'd754: row_of_pixels <= 8'b00000000;
		12'd755: row_of_pixels <= 8'b00000000;
		12'd756: row_of_pixels <= 8'b01000000;
		12'd757: row_of_pixels <= 8'b01100000;
		12'd758: row_of_pixels <= 8'b00110000;
		12'd759: row_of_pixels <= 8'b00011000;
		12'd760: row_of_pixels <= 8'b00001100;
		12'd761: row_of_pixels <= 8'b00000110;
		12'd762: row_of_pixels <= 8'b00000011;
		12'd763: row_of_pixels <= 8'b00000001;
		12'd764: row_of_pixels <= 8'b00000000;
		12'd765: row_of_pixels <= 8'b00000000;
		12'd766: row_of_pixels <= 8'b00000000;
		12'd767: row_of_pixels <= 8'b00000000;
		12'd768: row_of_pixels <= 8'b00000000;
		12'd769: row_of_pixels <= 8'b00000000;
		12'd770: row_of_pixels <= 8'b00111110;
		12'd771: row_of_pixels <= 8'b01100011;
		12'd772: row_of_pixels <= 8'b01100011;
		12'd773: row_of_pixels <= 8'b01110011;
		12'd774: row_of_pixels <= 8'b01111011;
		12'd775: row_of_pixels <= 8'b01101111;
		12'd776: row_of_pixels <= 8'b01100111;
		12'd777: row_of_pixels <= 8'b01100011;
		12'd778: row_of_pixels <= 8'b01100011;
		12'd779: row_of_pixels <= 8'b00111110;
		12'd780: row_of_pixels <= 8'b00000000;
		12'd781: row_of_pixels <= 8'b00000000;
		12'd782: row_of_pixels <= 8'b00000000;
		12'd783: row_of_pixels <= 8'b00000000;
		12'd784: row_of_pixels <= 8'b00000000;
		12'd785: row_of_pixels <= 8'b00000000;
		12'd786: row_of_pixels <= 8'b00011000;
		12'd787: row_of_pixels <= 8'b00011100;
		12'd788: row_of_pixels <= 8'b00011110;
		12'd789: row_of_pixels <= 8'b00011000;
		12'd790: row_of_pixels <= 8'b00011000;
		12'd791: row_of_pixels <= 8'b00011000;
		12'd792: row_of_pixels <= 8'b00011000;
		12'd793: row_of_pixels <= 8'b00011000;
		12'd794: row_of_pixels <= 8'b00011000;
		12'd795: row_of_pixels <= 8'b01111110;
		12'd796: row_of_pixels <= 8'b00000000;
		12'd797: row_of_pixels <= 8'b00000000;
		12'd798: row_of_pixels <= 8'b00000000;
		12'd799: row_of_pixels <= 8'b00000000;
		12'd800: row_of_pixels <= 8'b00000000;
		12'd801: row_of_pixels <= 8'b00000000;
		12'd802: row_of_pixels <= 8'b00111110;
		12'd803: row_of_pixels <= 8'b01100011;
		12'd804: row_of_pixels <= 8'b01100000;
		12'd805: row_of_pixels <= 8'b00110000;
		12'd806: row_of_pixels <= 8'b00011000;
		12'd807: row_of_pixels <= 8'b00001100;
		12'd808: row_of_pixels <= 8'b00000110;
		12'd809: row_of_pixels <= 8'b00000011;
		12'd810: row_of_pixels <= 8'b01100011;
		12'd811: row_of_pixels <= 8'b01111111;
		12'd812: row_of_pixels <= 8'b00000000;
		12'd813: row_of_pixels <= 8'b00000000;
		12'd814: row_of_pixels <= 8'b00000000;
		12'd815: row_of_pixels <= 8'b00000000;
		12'd816: row_of_pixels <= 8'b00000000;
		12'd817: row_of_pixels <= 8'b00000000;
		12'd818: row_of_pixels <= 8'b00111110;
		12'd819: row_of_pixels <= 8'b01100011;
		12'd820: row_of_pixels <= 8'b01100000;
		12'd821: row_of_pixels <= 8'b01100000;
		12'd822: row_of_pixels <= 8'b00111100;
		12'd823: row_of_pixels <= 8'b01100000;
		12'd824: row_of_pixels <= 8'b01100000;
		12'd825: row_of_pixels <= 8'b01100000;
		12'd826: row_of_pixels <= 8'b01100011;
		12'd827: row_of_pixels <= 8'b00111110;
		12'd828: row_of_pixels <= 8'b00000000;
		12'd829: row_of_pixels <= 8'b00000000;
		12'd830: row_of_pixels <= 8'b00000000;
		12'd831: row_of_pixels <= 8'b00000000;
		12'd832: row_of_pixels <= 8'b00000000;
		12'd833: row_of_pixels <= 8'b00000000;
		12'd834: row_of_pixels <= 8'b00110000;
		12'd835: row_of_pixels <= 8'b00111000;
		12'd836: row_of_pixels <= 8'b00111100;
		12'd837: row_of_pixels <= 8'b00110110;
		12'd838: row_of_pixels <= 8'b00110011;
		12'd839: row_of_pixels <= 8'b01111111;
		12'd840: row_of_pixels <= 8'b00110000;
		12'd841: row_of_pixels <= 8'b00110000;
		12'd842: row_of_pixels <= 8'b00110000;
		12'd843: row_of_pixels <= 8'b01111000;
		12'd844: row_of_pixels <= 8'b00000000;
		12'd845: row_of_pixels <= 8'b00000000;
		12'd846: row_of_pixels <= 8'b00000000;
		12'd847: row_of_pixels <= 8'b00000000;
		12'd848: row_of_pixels <= 8'b00000000;
		12'd849: row_of_pixels <= 8'b00000000;
		12'd850: row_of_pixels <= 8'b01111111;
		12'd851: row_of_pixels <= 8'b00000011;
		12'd852: row_of_pixels <= 8'b00000011;
		12'd853: row_of_pixels <= 8'b00000011;
		12'd854: row_of_pixels <= 8'b00111111;
		12'd855: row_of_pixels <= 8'b01100000;
		12'd856: row_of_pixels <= 8'b01100000;
		12'd857: row_of_pixels <= 8'b01100000;
		12'd858: row_of_pixels <= 8'b01100011;
		12'd859: row_of_pixels <= 8'b00111110;
		12'd860: row_of_pixels <= 8'b00000000;
		12'd861: row_of_pixels <= 8'b00000000;
		12'd862: row_of_pixels <= 8'b00000000;
		12'd863: row_of_pixels <= 8'b00000000;
		12'd864: row_of_pixels <= 8'b00000000;
		12'd865: row_of_pixels <= 8'b00000000;
		12'd866: row_of_pixels <= 8'b00011100;
		12'd867: row_of_pixels <= 8'b00000110;
		12'd868: row_of_pixels <= 8'b00000011;
		12'd869: row_of_pixels <= 8'b00000011;
		12'd870: row_of_pixels <= 8'b00111111;
		12'd871: row_of_pixels <= 8'b01100011;
		12'd872: row_of_pixels <= 8'b01100011;
		12'd873: row_of_pixels <= 8'b01100011;
		12'd874: row_of_pixels <= 8'b01100011;
		12'd875: row_of_pixels <= 8'b00111110;
		12'd876: row_of_pixels <= 8'b00000000;
		12'd877: row_of_pixels <= 8'b00000000;
		12'd878: row_of_pixels <= 8'b00000000;
		12'd879: row_of_pixels <= 8'b00000000;
		12'd880: row_of_pixels <= 8'b00000000;
		12'd881: row_of_pixels <= 8'b00000000;
		12'd882: row_of_pixels <= 8'b01111111;
		12'd883: row_of_pixels <= 8'b01100011;
		12'd884: row_of_pixels <= 8'b01100000;
		12'd885: row_of_pixels <= 8'b01100000;
		12'd886: row_of_pixels <= 8'b00110000;
		12'd887: row_of_pixels <= 8'b00011000;
		12'd888: row_of_pixels <= 8'b00001100;
		12'd889: row_of_pixels <= 8'b00001100;
		12'd890: row_of_pixels <= 8'b00001100;
		12'd891: row_of_pixels <= 8'b00001100;
		12'd892: row_of_pixels <= 8'b00000000;
		12'd893: row_of_pixels <= 8'b00000000;
		12'd894: row_of_pixels <= 8'b00000000;
		12'd895: row_of_pixels <= 8'b00000000;
		12'd896: row_of_pixels <= 8'b00000000;
		12'd897: row_of_pixels <= 8'b00000000;
		12'd898: row_of_pixels <= 8'b00111110;
		12'd899: row_of_pixels <= 8'b01100011;
		12'd900: row_of_pixels <= 8'b01100011;
		12'd901: row_of_pixels <= 8'b01100011;
		12'd902: row_of_pixels <= 8'b00111110;
		12'd903: row_of_pixels <= 8'b01100011;
		12'd904: row_of_pixels <= 8'b01100011;
		12'd905: row_of_pixels <= 8'b01100011;
		12'd906: row_of_pixels <= 8'b01100011;
		12'd907: row_of_pixels <= 8'b00111110;
		12'd908: row_of_pixels <= 8'b00000000;
		12'd909: row_of_pixels <= 8'b00000000;
		12'd910: row_of_pixels <= 8'b00000000;
		12'd911: row_of_pixels <= 8'b00000000;
		12'd912: row_of_pixels <= 8'b00000000;
		12'd913: row_of_pixels <= 8'b00000000;
		12'd914: row_of_pixels <= 8'b00111110;
		12'd915: row_of_pixels <= 8'b01100011;
		12'd916: row_of_pixels <= 8'b01100011;
		12'd917: row_of_pixels <= 8'b01100011;
		12'd918: row_of_pixels <= 8'b01111110;
		12'd919: row_of_pixels <= 8'b01100000;
		12'd920: row_of_pixels <= 8'b01100000;
		12'd921: row_of_pixels <= 8'b01100000;
		12'd922: row_of_pixels <= 8'b00110000;
		12'd923: row_of_pixels <= 8'b00011110;
		12'd924: row_of_pixels <= 8'b00000000;
		12'd925: row_of_pixels <= 8'b00000000;
		12'd926: row_of_pixels <= 8'b00000000;
		12'd927: row_of_pixels <= 8'b00000000;
		12'd928: row_of_pixels <= 8'b00000000;
		12'd929: row_of_pixels <= 8'b00000000;
		12'd930: row_of_pixels <= 8'b00000000;
		12'd931: row_of_pixels <= 8'b00000000;
		12'd932: row_of_pixels <= 8'b00011000;
		12'd933: row_of_pixels <= 8'b00011000;
		12'd934: row_of_pixels <= 8'b00000000;
		12'd935: row_of_pixels <= 8'b00000000;
		12'd936: row_of_pixels <= 8'b00000000;
		12'd937: row_of_pixels <= 8'b00011000;
		12'd938: row_of_pixels <= 8'b00011000;
		12'd939: row_of_pixels <= 8'b00000000;
		12'd940: row_of_pixels <= 8'b00000000;
		12'd941: row_of_pixels <= 8'b00000000;
		12'd942: row_of_pixels <= 8'b00000000;
		12'd943: row_of_pixels <= 8'b00000000;
		12'd944: row_of_pixels <= 8'b00000000;
		12'd945: row_of_pixels <= 8'b00000000;
		12'd946: row_of_pixels <= 8'b00000000;
		12'd947: row_of_pixels <= 8'b00000000;
		12'd948: row_of_pixels <= 8'b00011000;
		12'd949: row_of_pixels <= 8'b00011000;
		12'd950: row_of_pixels <= 8'b00000000;
		12'd951: row_of_pixels <= 8'b00000000;
		12'd952: row_of_pixels <= 8'b00000000;
		12'd953: row_of_pixels <= 8'b00011000;
		12'd954: row_of_pixels <= 8'b00011000;
		12'd955: row_of_pixels <= 8'b00001100;
		12'd956: row_of_pixels <= 8'b00000000;
		12'd957: row_of_pixels <= 8'b00000000;
		12'd958: row_of_pixels <= 8'b00000000;
		12'd959: row_of_pixels <= 8'b00000000;
		12'd960: row_of_pixels <= 8'b00000000;
		12'd961: row_of_pixels <= 8'b00000000;
		12'd962: row_of_pixels <= 8'b00000000;
		12'd963: row_of_pixels <= 8'b01100000;
		12'd964: row_of_pixels <= 8'b00110000;
		12'd965: row_of_pixels <= 8'b00011000;
		12'd966: row_of_pixels <= 8'b00001100;
		12'd967: row_of_pixels <= 8'b00000110;
		12'd968: row_of_pixels <= 8'b00001100;
		12'd969: row_of_pixels <= 8'b00011000;
		12'd970: row_of_pixels <= 8'b00110000;
		12'd971: row_of_pixels <= 8'b01100000;
		12'd972: row_of_pixels <= 8'b00000000;
		12'd973: row_of_pixels <= 8'b00000000;
		12'd974: row_of_pixels <= 8'b00000000;
		12'd975: row_of_pixels <= 8'b00000000;
		12'd976: row_of_pixels <= 8'b00000000;
		12'd977: row_of_pixels <= 8'b00000000;
		12'd978: row_of_pixels <= 8'b00000000;
		12'd979: row_of_pixels <= 8'b00000000;
		12'd980: row_of_pixels <= 8'b00000000;
		12'd981: row_of_pixels <= 8'b01111110;
		12'd982: row_of_pixels <= 8'b00000000;
		12'd983: row_of_pixels <= 8'b00000000;
		12'd984: row_of_pixels <= 8'b01111110;
		12'd985: row_of_pixels <= 8'b00000000;
		12'd986: row_of_pixels <= 8'b00000000;
		12'd987: row_of_pixels <= 8'b00000000;
		12'd988: row_of_pixels <= 8'b00000000;
		12'd989: row_of_pixels <= 8'b00000000;
		12'd990: row_of_pixels <= 8'b00000000;
		12'd991: row_of_pixels <= 8'b00000000;
		12'd992: row_of_pixels <= 8'b00000000;
		12'd993: row_of_pixels <= 8'b00000000;
		12'd994: row_of_pixels <= 8'b00000000;
		12'd995: row_of_pixels <= 8'b00000110;
		12'd996: row_of_pixels <= 8'b00001100;
		12'd997: row_of_pixels <= 8'b00011000;
		12'd998: row_of_pixels <= 8'b00110000;
		12'd999: row_of_pixels <= 8'b01100000;
		12'd1000: row_of_pixels <= 8'b00110000;
		12'd1001: row_of_pixels <= 8'b00011000;
		12'd1002: row_of_pixels <= 8'b00001100;
		12'd1003: row_of_pixels <= 8'b00000110;
		12'd1004: row_of_pixels <= 8'b00000000;
		12'd1005: row_of_pixels <= 8'b00000000;
		12'd1006: row_of_pixels <= 8'b00000000;
		12'd1007: row_of_pixels <= 8'b00000000;
		12'd1008: row_of_pixels <= 8'b00000000;
		12'd1009: row_of_pixels <= 8'b00000000;
		12'd1010: row_of_pixels <= 8'b00111110;
		12'd1011: row_of_pixels <= 8'b01100011;
		12'd1012: row_of_pixels <= 8'b01100011;
		12'd1013: row_of_pixels <= 8'b00110000;
		12'd1014: row_of_pixels <= 8'b00011000;
		12'd1015: row_of_pixels <= 8'b00011000;
		12'd1016: row_of_pixels <= 8'b00011000;
		12'd1017: row_of_pixels <= 8'b00000000;
		12'd1018: row_of_pixels <= 8'b00011000;
		12'd1019: row_of_pixels <= 8'b00011000;
		12'd1020: row_of_pixels <= 8'b00000000;
		12'd1021: row_of_pixels <= 8'b00000000;
		12'd1022: row_of_pixels <= 8'b00000000;
		12'd1023: row_of_pixels <= 8'b00000000;
		12'd1024: row_of_pixels <= 8'b00000000;
		12'd1025: row_of_pixels <= 8'b00000000;
		12'd1026: row_of_pixels <= 8'b00111110;
		12'd1027: row_of_pixels <= 8'b01100011;
		12'd1028: row_of_pixels <= 8'b01100011;
		12'd1029: row_of_pixels <= 8'b01100011;
		12'd1030: row_of_pixels <= 8'b01111011;
		12'd1031: row_of_pixels <= 8'b01111011;
		12'd1032: row_of_pixels <= 8'b01111011;
		12'd1033: row_of_pixels <= 8'b00111011;
		12'd1034: row_of_pixels <= 8'b00000011;
		12'd1035: row_of_pixels <= 8'b00111110;
		12'd1036: row_of_pixels <= 8'b00000000;
		12'd1037: row_of_pixels <= 8'b00000000;
		12'd1038: row_of_pixels <= 8'b00000000;
		12'd1039: row_of_pixels <= 8'b00000000;
		12'd1040: row_of_pixels <= 8'b00000000;
		12'd1041: row_of_pixels <= 8'b00000000;
		12'd1042: row_of_pixels <= 8'b00001000;
		12'd1043: row_of_pixels <= 8'b00011100;
		12'd1044: row_of_pixels <= 8'b00110110;
		12'd1045: row_of_pixels <= 8'b01100011;
		12'd1046: row_of_pixels <= 8'b01100011;
		12'd1047: row_of_pixels <= 8'b01111111;
		12'd1048: row_of_pixels <= 8'b01100011;
		12'd1049: row_of_pixels <= 8'b01100011;
		12'd1050: row_of_pixels <= 8'b01100011;
		12'd1051: row_of_pixels <= 8'b01100011;
		12'd1052: row_of_pixels <= 8'b00000000;
		12'd1053: row_of_pixels <= 8'b00000000;
		12'd1054: row_of_pixels <= 8'b00000000;
		12'd1055: row_of_pixels <= 8'b00000000;
		12'd1056: row_of_pixels <= 8'b00000000;
		12'd1057: row_of_pixels <= 8'b00000000;
		12'd1058: row_of_pixels <= 8'b00111111;
		12'd1059: row_of_pixels <= 8'b01100110;
		12'd1060: row_of_pixels <= 8'b01100110;
		12'd1061: row_of_pixels <= 8'b01100110;
		12'd1062: row_of_pixels <= 8'b00111110;
		12'd1063: row_of_pixels <= 8'b01100110;
		12'd1064: row_of_pixels <= 8'b01100110;
		12'd1065: row_of_pixels <= 8'b01100110;
		12'd1066: row_of_pixels <= 8'b01100110;
		12'd1067: row_of_pixels <= 8'b00111111;
		12'd1068: row_of_pixels <= 8'b00000000;
		12'd1069: row_of_pixels <= 8'b00000000;
		12'd1070: row_of_pixels <= 8'b00000000;
		12'd1071: row_of_pixels <= 8'b00000000;
		12'd1072: row_of_pixels <= 8'b00000000;
		12'd1073: row_of_pixels <= 8'b00000000;
		12'd1074: row_of_pixels <= 8'b00111100;
		12'd1075: row_of_pixels <= 8'b01100110;
		12'd1076: row_of_pixels <= 8'b01000011;
		12'd1077: row_of_pixels <= 8'b00000011;
		12'd1078: row_of_pixels <= 8'b00000011;
		12'd1079: row_of_pixels <= 8'b00000011;
		12'd1080: row_of_pixels <= 8'b00000011;
		12'd1081: row_of_pixels <= 8'b01000011;
		12'd1082: row_of_pixels <= 8'b01100110;
		12'd1083: row_of_pixels <= 8'b00111100;
		12'd1084: row_of_pixels <= 8'b00000000;
		12'd1085: row_of_pixels <= 8'b00000000;
		12'd1086: row_of_pixels <= 8'b00000000;
		12'd1087: row_of_pixels <= 8'b00000000;
		12'd1088: row_of_pixels <= 8'b00000000;
		12'd1089: row_of_pixels <= 8'b00000000;
		12'd1090: row_of_pixels <= 8'b00011111;
		12'd1091: row_of_pixels <= 8'b00110110;
		12'd1092: row_of_pixels <= 8'b01100110;
		12'd1093: row_of_pixels <= 8'b01100110;
		12'd1094: row_of_pixels <= 8'b01100110;
		12'd1095: row_of_pixels <= 8'b01100110;
		12'd1096: row_of_pixels <= 8'b01100110;
		12'd1097: row_of_pixels <= 8'b01100110;
		12'd1098: row_of_pixels <= 8'b00110110;
		12'd1099: row_of_pixels <= 8'b00011111;
		12'd1100: row_of_pixels <= 8'b00000000;
		12'd1101: row_of_pixels <= 8'b00000000;
		12'd1102: row_of_pixels <= 8'b00000000;
		12'd1103: row_of_pixels <= 8'b00000000;
		12'd1104: row_of_pixels <= 8'b00000000;
		12'd1105: row_of_pixels <= 8'b00000000;
		12'd1106: row_of_pixels <= 8'b01111111;
		12'd1107: row_of_pixels <= 8'b01100110;
		12'd1108: row_of_pixels <= 8'b01000110;
		12'd1109: row_of_pixels <= 8'b00010110;
		12'd1110: row_of_pixels <= 8'b00011110;
		12'd1111: row_of_pixels <= 8'b00010110;
		12'd1112: row_of_pixels <= 8'b00000110;
		12'd1113: row_of_pixels <= 8'b01000110;
		12'd1114: row_of_pixels <= 8'b01100110;
		12'd1115: row_of_pixels <= 8'b01111111;
		12'd1116: row_of_pixels <= 8'b00000000;
		12'd1117: row_of_pixels <= 8'b00000000;
		12'd1118: row_of_pixels <= 8'b00000000;
		12'd1119: row_of_pixels <= 8'b00000000;
		12'd1120: row_of_pixels <= 8'b00000000;
		12'd1121: row_of_pixels <= 8'b00000000;
		12'd1122: row_of_pixels <= 8'b01111111;
		12'd1123: row_of_pixels <= 8'b01100110;
		12'd1124: row_of_pixels <= 8'b01000110;
		12'd1125: row_of_pixels <= 8'b00010110;
		12'd1126: row_of_pixels <= 8'b00011110;
		12'd1127: row_of_pixels <= 8'b00010110;
		12'd1128: row_of_pixels <= 8'b00000110;
		12'd1129: row_of_pixels <= 8'b00000110;
		12'd1130: row_of_pixels <= 8'b00000110;
		12'd1131: row_of_pixels <= 8'b00001111;
		12'd1132: row_of_pixels <= 8'b00000000;
		12'd1133: row_of_pixels <= 8'b00000000;
		12'd1134: row_of_pixels <= 8'b00000000;
		12'd1135: row_of_pixels <= 8'b00000000;
		12'd1136: row_of_pixels <= 8'b00000000;
		12'd1137: row_of_pixels <= 8'b00000000;
		12'd1138: row_of_pixels <= 8'b00111100;
		12'd1139: row_of_pixels <= 8'b01100110;
		12'd1140: row_of_pixels <= 8'b01000011;
		12'd1141: row_of_pixels <= 8'b00000011;
		12'd1142: row_of_pixels <= 8'b00000011;
		12'd1143: row_of_pixels <= 8'b01111011;
		12'd1144: row_of_pixels <= 8'b01100011;
		12'd1145: row_of_pixels <= 8'b01100011;
		12'd1146: row_of_pixels <= 8'b01100110;
		12'd1147: row_of_pixels <= 8'b01011100;
		12'd1148: row_of_pixels <= 8'b00000000;
		12'd1149: row_of_pixels <= 8'b00000000;
		12'd1150: row_of_pixels <= 8'b00000000;
		12'd1151: row_of_pixels <= 8'b00000000;
		12'd1152: row_of_pixels <= 8'b00000000;
		12'd1153: row_of_pixels <= 8'b00000000;
		12'd1154: row_of_pixels <= 8'b01100011;
		12'd1155: row_of_pixels <= 8'b01100011;
		12'd1156: row_of_pixels <= 8'b01100011;
		12'd1157: row_of_pixels <= 8'b01100011;
		12'd1158: row_of_pixels <= 8'b01111111;
		12'd1159: row_of_pixels <= 8'b01100011;
		12'd1160: row_of_pixels <= 8'b01100011;
		12'd1161: row_of_pixels <= 8'b01100011;
		12'd1162: row_of_pixels <= 8'b01100011;
		12'd1163: row_of_pixels <= 8'b01100011;
		12'd1164: row_of_pixels <= 8'b00000000;
		12'd1165: row_of_pixels <= 8'b00000000;
		12'd1166: row_of_pixels <= 8'b00000000;
		12'd1167: row_of_pixels <= 8'b00000000;
		12'd1168: row_of_pixels <= 8'b00000000;
		12'd1169: row_of_pixels <= 8'b00000000;
		12'd1170: row_of_pixels <= 8'b00111100;
		12'd1171: row_of_pixels <= 8'b00011000;
		12'd1172: row_of_pixels <= 8'b00011000;
		12'd1173: row_of_pixels <= 8'b00011000;
		12'd1174: row_of_pixels <= 8'b00011000;
		12'd1175: row_of_pixels <= 8'b00011000;
		12'd1176: row_of_pixels <= 8'b00011000;
		12'd1177: row_of_pixels <= 8'b00011000;
		12'd1178: row_of_pixels <= 8'b00011000;
		12'd1179: row_of_pixels <= 8'b00111100;
		12'd1180: row_of_pixels <= 8'b00000000;
		12'd1181: row_of_pixels <= 8'b00000000;
		12'd1182: row_of_pixels <= 8'b00000000;
		12'd1183: row_of_pixels <= 8'b00000000;
		12'd1184: row_of_pixels <= 8'b00000000;
		12'd1185: row_of_pixels <= 8'b00000000;
		12'd1186: row_of_pixels <= 8'b01111000;
		12'd1187: row_of_pixels <= 8'b00110000;
		12'd1188: row_of_pixels <= 8'b00110000;
		12'd1189: row_of_pixels <= 8'b00110000;
		12'd1190: row_of_pixels <= 8'b00110000;
		12'd1191: row_of_pixels <= 8'b00110000;
		12'd1192: row_of_pixels <= 8'b00110011;
		12'd1193: row_of_pixels <= 8'b00110011;
		12'd1194: row_of_pixels <= 8'b00110011;
		12'd1195: row_of_pixels <= 8'b00011110;
		12'd1196: row_of_pixels <= 8'b00000000;
		12'd1197: row_of_pixels <= 8'b00000000;
		12'd1198: row_of_pixels <= 8'b00000000;
		12'd1199: row_of_pixels <= 8'b00000000;
		12'd1200: row_of_pixels <= 8'b00000000;
		12'd1201: row_of_pixels <= 8'b00000000;
		12'd1202: row_of_pixels <= 8'b01100111;
		12'd1203: row_of_pixels <= 8'b01100110;
		12'd1204: row_of_pixels <= 8'b01100110;
		12'd1205: row_of_pixels <= 8'b00110110;
		12'd1206: row_of_pixels <= 8'b00011110;
		12'd1207: row_of_pixels <= 8'b00011110;
		12'd1208: row_of_pixels <= 8'b00110110;
		12'd1209: row_of_pixels <= 8'b01100110;
		12'd1210: row_of_pixels <= 8'b01100110;
		12'd1211: row_of_pixels <= 8'b01100111;
		12'd1212: row_of_pixels <= 8'b00000000;
		12'd1213: row_of_pixels <= 8'b00000000;
		12'd1214: row_of_pixels <= 8'b00000000;
		12'd1215: row_of_pixels <= 8'b00000000;
		12'd1216: row_of_pixels <= 8'b00000000;
		12'd1217: row_of_pixels <= 8'b00000000;
		12'd1218: row_of_pixels <= 8'b00001111;
		12'd1219: row_of_pixels <= 8'b00000110;
		12'd1220: row_of_pixels <= 8'b00000110;
		12'd1221: row_of_pixels <= 8'b00000110;
		12'd1222: row_of_pixels <= 8'b00000110;
		12'd1223: row_of_pixels <= 8'b00000110;
		12'd1224: row_of_pixels <= 8'b00000110;
		12'd1225: row_of_pixels <= 8'b01000110;
		12'd1226: row_of_pixels <= 8'b01100110;
		12'd1227: row_of_pixels <= 8'b01111111;
		12'd1228: row_of_pixels <= 8'b00000000;
		12'd1229: row_of_pixels <= 8'b00000000;
		12'd1230: row_of_pixels <= 8'b00000000;
		12'd1231: row_of_pixels <= 8'b00000000;
		12'd1232: row_of_pixels <= 8'b00000000;
		12'd1233: row_of_pixels <= 8'b00000000;
		12'd1234: row_of_pixels <= 8'b11000011;
		12'd1235: row_of_pixels <= 8'b11100111;
		12'd1236: row_of_pixels <= 8'b11111111;
		12'd1237: row_of_pixels <= 8'b11111111;
		12'd1238: row_of_pixels <= 8'b11011011;
		12'd1239: row_of_pixels <= 8'b11000011;
		12'd1240: row_of_pixels <= 8'b11000011;
		12'd1241: row_of_pixels <= 8'b11000011;
		12'd1242: row_of_pixels <= 8'b11000011;
		12'd1243: row_of_pixels <= 8'b11000011;
		12'd1244: row_of_pixels <= 8'b00000000;
		12'd1245: row_of_pixels <= 8'b00000000;
		12'd1246: row_of_pixels <= 8'b00000000;
		12'd1247: row_of_pixels <= 8'b00000000;
		12'd1248: row_of_pixels <= 8'b00000000;
		12'd1249: row_of_pixels <= 8'b00000000;
		12'd1250: row_of_pixels <= 8'b01100011;
		12'd1251: row_of_pixels <= 8'b01100111;
		12'd1252: row_of_pixels <= 8'b01101111;
		12'd1253: row_of_pixels <= 8'b01111111;
		12'd1254: row_of_pixels <= 8'b01111011;
		12'd1255: row_of_pixels <= 8'b01110011;
		12'd1256: row_of_pixels <= 8'b01100011;
		12'd1257: row_of_pixels <= 8'b01100011;
		12'd1258: row_of_pixels <= 8'b01100011;
		12'd1259: row_of_pixels <= 8'b01100011;
		12'd1260: row_of_pixels <= 8'b00000000;
		12'd1261: row_of_pixels <= 8'b00000000;
		12'd1262: row_of_pixels <= 8'b00000000;
		12'd1263: row_of_pixels <= 8'b00000000;
		12'd1264: row_of_pixels <= 8'b00000000;
		12'd1265: row_of_pixels <= 8'b00000000;
		12'd1266: row_of_pixels <= 8'b00111110;
		12'd1267: row_of_pixels <= 8'b01100011;
		12'd1268: row_of_pixels <= 8'b01100011;
		12'd1269: row_of_pixels <= 8'b01100011;
		12'd1270: row_of_pixels <= 8'b01100011;
		12'd1271: row_of_pixels <= 8'b01100011;
		12'd1272: row_of_pixels <= 8'b01100011;
		12'd1273: row_of_pixels <= 8'b01100011;
		12'd1274: row_of_pixels <= 8'b01100011;
		12'd1275: row_of_pixels <= 8'b00111110;
		12'd1276: row_of_pixels <= 8'b00000000;
		12'd1277: row_of_pixels <= 8'b00000000;
		12'd1278: row_of_pixels <= 8'b00000000;
		12'd1279: row_of_pixels <= 8'b00000000;
		12'd1280: row_of_pixels <= 8'b00000000;
		12'd1281: row_of_pixels <= 8'b00000000;
		12'd1282: row_of_pixels <= 8'b00111111;
		12'd1283: row_of_pixels <= 8'b01100110;
		12'd1284: row_of_pixels <= 8'b01100110;
		12'd1285: row_of_pixels <= 8'b01100110;
		12'd1286: row_of_pixels <= 8'b00111110;
		12'd1287: row_of_pixels <= 8'b00000110;
		12'd1288: row_of_pixels <= 8'b00000110;
		12'd1289: row_of_pixels <= 8'b00000110;
		12'd1290: row_of_pixels <= 8'b00000110;
		12'd1291: row_of_pixels <= 8'b00001111;
		12'd1292: row_of_pixels <= 8'b00000000;
		12'd1293: row_of_pixels <= 8'b00000000;
		12'd1294: row_of_pixels <= 8'b00000000;
		12'd1295: row_of_pixels <= 8'b00000000;
		12'd1296: row_of_pixels <= 8'b00000000;
		12'd1297: row_of_pixels <= 8'b00000000;
		12'd1298: row_of_pixels <= 8'b00111110;
		12'd1299: row_of_pixels <= 8'b01100011;
		12'd1300: row_of_pixels <= 8'b01100011;
		12'd1301: row_of_pixels <= 8'b01100011;
		12'd1302: row_of_pixels <= 8'b01100011;
		12'd1303: row_of_pixels <= 8'b01100011;
		12'd1304: row_of_pixels <= 8'b01100011;
		12'd1305: row_of_pixels <= 8'b01101011;
		12'd1306: row_of_pixels <= 8'b01111011;
		12'd1307: row_of_pixels <= 8'b00111110;
		12'd1308: row_of_pixels <= 8'b00110000;
		12'd1309: row_of_pixels <= 8'b01110000;
		12'd1310: row_of_pixels <= 8'b00000000;
		12'd1311: row_of_pixels <= 8'b00000000;
		12'd1312: row_of_pixels <= 8'b00000000;
		12'd1313: row_of_pixels <= 8'b00000000;
		12'd1314: row_of_pixels <= 8'b00111111;
		12'd1315: row_of_pixels <= 8'b01100110;
		12'd1316: row_of_pixels <= 8'b01100110;
		12'd1317: row_of_pixels <= 8'b01100110;
		12'd1318: row_of_pixels <= 8'b00111110;
		12'd1319: row_of_pixels <= 8'b00110110;
		12'd1320: row_of_pixels <= 8'b01100110;
		12'd1321: row_of_pixels <= 8'b01100110;
		12'd1322: row_of_pixels <= 8'b01100110;
		12'd1323: row_of_pixels <= 8'b01100111;
		12'd1324: row_of_pixels <= 8'b00000000;
		12'd1325: row_of_pixels <= 8'b00000000;
		12'd1326: row_of_pixels <= 8'b00000000;
		12'd1327: row_of_pixels <= 8'b00000000;
		12'd1328: row_of_pixels <= 8'b00000000;
		12'd1329: row_of_pixels <= 8'b00000000;
		12'd1330: row_of_pixels <= 8'b00111110;
		12'd1331: row_of_pixels <= 8'b01100011;
		12'd1332: row_of_pixels <= 8'b01100011;
		12'd1333: row_of_pixels <= 8'b00000110;
		12'd1334: row_of_pixels <= 8'b00011100;
		12'd1335: row_of_pixels <= 8'b00110000;
		12'd1336: row_of_pixels <= 8'b01100000;
		12'd1337: row_of_pixels <= 8'b01100011;
		12'd1338: row_of_pixels <= 8'b01100011;
		12'd1339: row_of_pixels <= 8'b00111110;
		12'd1340: row_of_pixels <= 8'b00000000;
		12'd1341: row_of_pixels <= 8'b00000000;
		12'd1342: row_of_pixels <= 8'b00000000;
		12'd1343: row_of_pixels <= 8'b00000000;
		12'd1344: row_of_pixels <= 8'b00000000;
		12'd1345: row_of_pixels <= 8'b00000000;
		12'd1346: row_of_pixels <= 8'b11111111;
		12'd1347: row_of_pixels <= 8'b11011011;
		12'd1348: row_of_pixels <= 8'b10011001;
		12'd1349: row_of_pixels <= 8'b00011000;
		12'd1350: row_of_pixels <= 8'b00011000;
		12'd1351: row_of_pixels <= 8'b00011000;
		12'd1352: row_of_pixels <= 8'b00011000;
		12'd1353: row_of_pixels <= 8'b00011000;
		12'd1354: row_of_pixels <= 8'b00011000;
		12'd1355: row_of_pixels <= 8'b00111100;
		12'd1356: row_of_pixels <= 8'b00000000;
		12'd1357: row_of_pixels <= 8'b00000000;
		12'd1358: row_of_pixels <= 8'b00000000;
		12'd1359: row_of_pixels <= 8'b00000000;
		12'd1360: row_of_pixels <= 8'b00000000;
		12'd1361: row_of_pixels <= 8'b00000000;
		12'd1362: row_of_pixels <= 8'b01100011;
		12'd1363: row_of_pixels <= 8'b01100011;
		12'd1364: row_of_pixels <= 8'b01100011;
		12'd1365: row_of_pixels <= 8'b01100011;
		12'd1366: row_of_pixels <= 8'b01100011;
		12'd1367: row_of_pixels <= 8'b01100011;
		12'd1368: row_of_pixels <= 8'b01100011;
		12'd1369: row_of_pixels <= 8'b01100011;
		12'd1370: row_of_pixels <= 8'b01100011;
		12'd1371: row_of_pixels <= 8'b00111110;
		12'd1372: row_of_pixels <= 8'b00000000;
		12'd1373: row_of_pixels <= 8'b00000000;
		12'd1374: row_of_pixels <= 8'b00000000;
		12'd1375: row_of_pixels <= 8'b00000000;
		12'd1376: row_of_pixels <= 8'b00000000;
		12'd1377: row_of_pixels <= 8'b00000000;
		12'd1378: row_of_pixels <= 8'b11000011;
		12'd1379: row_of_pixels <= 8'b11000011;
		12'd1380: row_of_pixels <= 8'b11000011;
		12'd1381: row_of_pixels <= 8'b11000011;
		12'd1382: row_of_pixels <= 8'b11000011;
		12'd1383: row_of_pixels <= 8'b11000011;
		12'd1384: row_of_pixels <= 8'b11000011;
		12'd1385: row_of_pixels <= 8'b01100110;
		12'd1386: row_of_pixels <= 8'b00111100;
		12'd1387: row_of_pixels <= 8'b00011000;
		12'd1388: row_of_pixels <= 8'b00000000;
		12'd1389: row_of_pixels <= 8'b00000000;
		12'd1390: row_of_pixels <= 8'b00000000;
		12'd1391: row_of_pixels <= 8'b00000000;
		12'd1392: row_of_pixels <= 8'b00000000;
		12'd1393: row_of_pixels <= 8'b00000000;
		12'd1394: row_of_pixels <= 8'b11000011;
		12'd1395: row_of_pixels <= 8'b11000011;
		12'd1396: row_of_pixels <= 8'b11000011;
		12'd1397: row_of_pixels <= 8'b11000011;
		12'd1398: row_of_pixels <= 8'b11000011;
		12'd1399: row_of_pixels <= 8'b11011011;
		12'd1400: row_of_pixels <= 8'b11011011;
		12'd1401: row_of_pixels <= 8'b11111111;
		12'd1402: row_of_pixels <= 8'b01100110;
		12'd1403: row_of_pixels <= 8'b01100110;
		12'd1404: row_of_pixels <= 8'b00000000;
		12'd1405: row_of_pixels <= 8'b00000000;
		12'd1406: row_of_pixels <= 8'b00000000;
		12'd1407: row_of_pixels <= 8'b00000000;
		12'd1408: row_of_pixels <= 8'b00000000;
		12'd1409: row_of_pixels <= 8'b00000000;
		12'd1410: row_of_pixels <= 8'b11000011;
		12'd1411: row_of_pixels <= 8'b11000011;
		12'd1412: row_of_pixels <= 8'b01100110;
		12'd1413: row_of_pixels <= 8'b00111100;
		12'd1414: row_of_pixels <= 8'b00011000;
		12'd1415: row_of_pixels <= 8'b00011000;
		12'd1416: row_of_pixels <= 8'b00111100;
		12'd1417: row_of_pixels <= 8'b01100110;
		12'd1418: row_of_pixels <= 8'b11000011;
		12'd1419: row_of_pixels <= 8'b11000011;
		12'd1420: row_of_pixels <= 8'b00000000;
		12'd1421: row_of_pixels <= 8'b00000000;
		12'd1422: row_of_pixels <= 8'b00000000;
		12'd1423: row_of_pixels <= 8'b00000000;
		12'd1424: row_of_pixels <= 8'b00000000;
		12'd1425: row_of_pixels <= 8'b00000000;
		12'd1426: row_of_pixels <= 8'b11000011;
		12'd1427: row_of_pixels <= 8'b11000011;
		12'd1428: row_of_pixels <= 8'b11000011;
		12'd1429: row_of_pixels <= 8'b01100110;
		12'd1430: row_of_pixels <= 8'b00111100;
		12'd1431: row_of_pixels <= 8'b00011000;
		12'd1432: row_of_pixels <= 8'b00011000;
		12'd1433: row_of_pixels <= 8'b00011000;
		12'd1434: row_of_pixels <= 8'b00011000;
		12'd1435: row_of_pixels <= 8'b00111100;
		12'd1436: row_of_pixels <= 8'b00000000;
		12'd1437: row_of_pixels <= 8'b00000000;
		12'd1438: row_of_pixels <= 8'b00000000;
		12'd1439: row_of_pixels <= 8'b00000000;
		12'd1440: row_of_pixels <= 8'b00000000;
		12'd1441: row_of_pixels <= 8'b00000000;
		12'd1442: row_of_pixels <= 8'b11111111;
		12'd1443: row_of_pixels <= 8'b11000011;
		12'd1444: row_of_pixels <= 8'b01100001;
		12'd1445: row_of_pixels <= 8'b00110000;
		12'd1446: row_of_pixels <= 8'b00011000;
		12'd1447: row_of_pixels <= 8'b00001100;
		12'd1448: row_of_pixels <= 8'b00000110;
		12'd1449: row_of_pixels <= 8'b10000011;
		12'd1450: row_of_pixels <= 8'b11000011;
		12'd1451: row_of_pixels <= 8'b11111111;
		12'd1452: row_of_pixels <= 8'b00000000;
		12'd1453: row_of_pixels <= 8'b00000000;
		12'd1454: row_of_pixels <= 8'b00000000;
		12'd1455: row_of_pixels <= 8'b00000000;
		12'd1456: row_of_pixels <= 8'b00000000;
		12'd1457: row_of_pixels <= 8'b00000000;
		12'd1458: row_of_pixels <= 8'b00111100;
		12'd1459: row_of_pixels <= 8'b00001100;
		12'd1460: row_of_pixels <= 8'b00001100;
		12'd1461: row_of_pixels <= 8'b00001100;
		12'd1462: row_of_pixels <= 8'b00001100;
		12'd1463: row_of_pixels <= 8'b00001100;
		12'd1464: row_of_pixels <= 8'b00001100;
		12'd1465: row_of_pixels <= 8'b00001100;
		12'd1466: row_of_pixels <= 8'b00001100;
		12'd1467: row_of_pixels <= 8'b00111100;
		12'd1468: row_of_pixels <= 8'b00000000;
		12'd1469: row_of_pixels <= 8'b00000000;
		12'd1470: row_of_pixels <= 8'b00000000;
		12'd1471: row_of_pixels <= 8'b00000000;
		12'd1472: row_of_pixels <= 8'b00000000;
		12'd1473: row_of_pixels <= 8'b00000000;
		12'd1474: row_of_pixels <= 8'b00000000;
		12'd1475: row_of_pixels <= 8'b00000001;
		12'd1476: row_of_pixels <= 8'b00000011;
		12'd1477: row_of_pixels <= 8'b00000111;
		12'd1478: row_of_pixels <= 8'b00001110;
		12'd1479: row_of_pixels <= 8'b00011100;
		12'd1480: row_of_pixels <= 8'b00111000;
		12'd1481: row_of_pixels <= 8'b01110000;
		12'd1482: row_of_pixels <= 8'b01100000;
		12'd1483: row_of_pixels <= 8'b01000000;
		12'd1484: row_of_pixels <= 8'b00000000;
		12'd1485: row_of_pixels <= 8'b00000000;
		12'd1486: row_of_pixels <= 8'b00000000;
		12'd1487: row_of_pixels <= 8'b00000000;
		12'd1488: row_of_pixels <= 8'b00000000;
		12'd1489: row_of_pixels <= 8'b00000000;
		12'd1490: row_of_pixels <= 8'b00111100;
		12'd1491: row_of_pixels <= 8'b00110000;
		12'd1492: row_of_pixels <= 8'b00110000;
		12'd1493: row_of_pixels <= 8'b00110000;
		12'd1494: row_of_pixels <= 8'b00110000;
		12'd1495: row_of_pixels <= 8'b00110000;
		12'd1496: row_of_pixels <= 8'b00110000;
		12'd1497: row_of_pixels <= 8'b00110000;
		12'd1498: row_of_pixels <= 8'b00110000;
		12'd1499: row_of_pixels <= 8'b00111100;
		12'd1500: row_of_pixels <= 8'b00000000;
		12'd1501: row_of_pixels <= 8'b00000000;
		12'd1502: row_of_pixels <= 8'b00000000;
		12'd1503: row_of_pixels <= 8'b00000000;
		12'd1504: row_of_pixels <= 8'b00001000;
		12'd1505: row_of_pixels <= 8'b00011100;
		12'd1506: row_of_pixels <= 8'b00110110;
		12'd1507: row_of_pixels <= 8'b01100011;
		12'd1508: row_of_pixels <= 8'b00000000;
		12'd1509: row_of_pixels <= 8'b00000000;
		12'd1510: row_of_pixels <= 8'b00000000;
		12'd1511: row_of_pixels <= 8'b00000000;
		12'd1512: row_of_pixels <= 8'b00000000;
		12'd1513: row_of_pixels <= 8'b00000000;
		12'd1514: row_of_pixels <= 8'b00000000;
		12'd1515: row_of_pixels <= 8'b00000000;
		12'd1516: row_of_pixels <= 8'b00000000;
		12'd1517: row_of_pixels <= 8'b00000000;
		12'd1518: row_of_pixels <= 8'b00000000;
		12'd1519: row_of_pixels <= 8'b00000000;
		12'd1520: row_of_pixels <= 8'b00000000;
		12'd1521: row_of_pixels <= 8'b00000000;
		12'd1522: row_of_pixels <= 8'b00000000;
		12'd1523: row_of_pixels <= 8'b00000000;
		12'd1524: row_of_pixels <= 8'b00000000;
		12'd1525: row_of_pixels <= 8'b00000000;
		12'd1526: row_of_pixels <= 8'b00000000;
		12'd1527: row_of_pixels <= 8'b00000000;
		12'd1528: row_of_pixels <= 8'b00000000;
		12'd1529: row_of_pixels <= 8'b00000000;
		12'd1530: row_of_pixels <= 8'b00000000;
		12'd1531: row_of_pixels <= 8'b00000000;
		12'd1532: row_of_pixels <= 8'b00000000;
		12'd1533: row_of_pixels <= 8'b11111111;
		12'd1534: row_of_pixels <= 8'b00000000;
		12'd1535: row_of_pixels <= 8'b00000000;
		12'd1536: row_of_pixels <= 8'b00001100;
		12'd1537: row_of_pixels <= 8'b00001100;
		12'd1538: row_of_pixels <= 8'b00011000;
		12'd1539: row_of_pixels <= 8'b00000000;
		12'd1540: row_of_pixels <= 8'b00000000;
		12'd1541: row_of_pixels <= 8'b00000000;
		12'd1542: row_of_pixels <= 8'b00000000;
		12'd1543: row_of_pixels <= 8'b00000000;
		12'd1544: row_of_pixels <= 8'b00000000;
		12'd1545: row_of_pixels <= 8'b00000000;
		12'd1546: row_of_pixels <= 8'b00000000;
		12'd1547: row_of_pixels <= 8'b00000000;
		12'd1548: row_of_pixels <= 8'b00000000;
		12'd1549: row_of_pixels <= 8'b00000000;
		12'd1550: row_of_pixels <= 8'b00000000;
		12'd1551: row_of_pixels <= 8'b00000000;
		12'd1552: row_of_pixels <= 8'b00000000;
		12'd1553: row_of_pixels <= 8'b00000000;
		12'd1554: row_of_pixels <= 8'b00000000;
		12'd1555: row_of_pixels <= 8'b00000000;
		12'd1556: row_of_pixels <= 8'b00000000;
		12'd1557: row_of_pixels <= 8'b00011110;
		12'd1558: row_of_pixels <= 8'b00110000;
		12'd1559: row_of_pixels <= 8'b00111110;
		12'd1560: row_of_pixels <= 8'b00110011;
		12'd1561: row_of_pixels <= 8'b00110011;
		12'd1562: row_of_pixels <= 8'b00110011;
		12'd1563: row_of_pixels <= 8'b01101110;
		12'd1564: row_of_pixels <= 8'b00000000;
		12'd1565: row_of_pixels <= 8'b00000000;
		12'd1566: row_of_pixels <= 8'b00000000;
		12'd1567: row_of_pixels <= 8'b00000000;
		12'd1568: row_of_pixels <= 8'b00000000;
		12'd1569: row_of_pixels <= 8'b00000000;
		12'd1570: row_of_pixels <= 8'b00000111;
		12'd1571: row_of_pixels <= 8'b00000110;
		12'd1572: row_of_pixels <= 8'b00000110;
		12'd1573: row_of_pixels <= 8'b00011110;
		12'd1574: row_of_pixels <= 8'b00110110;
		12'd1575: row_of_pixels <= 8'b01100110;
		12'd1576: row_of_pixels <= 8'b01100110;
		12'd1577: row_of_pixels <= 8'b01100110;
		12'd1578: row_of_pixels <= 8'b01100110;
		12'd1579: row_of_pixels <= 8'b00111110;
		12'd1580: row_of_pixels <= 8'b00000000;
		12'd1581: row_of_pixels <= 8'b00000000;
		12'd1582: row_of_pixels <= 8'b00000000;
		12'd1583: row_of_pixels <= 8'b00000000;
		12'd1584: row_of_pixels <= 8'b00000000;
		12'd1585: row_of_pixels <= 8'b00000000;
		12'd1586: row_of_pixels <= 8'b00000000;
		12'd1587: row_of_pixels <= 8'b00000000;
		12'd1588: row_of_pixels <= 8'b00000000;
		12'd1589: row_of_pixels <= 8'b00111110;
		12'd1590: row_of_pixels <= 8'b01100011;
		12'd1591: row_of_pixels <= 8'b00000011;
		12'd1592: row_of_pixels <= 8'b00000011;
		12'd1593: row_of_pixels <= 8'b00000011;
		12'd1594: row_of_pixels <= 8'b01100011;
		12'd1595: row_of_pixels <= 8'b00111110;
		12'd1596: row_of_pixels <= 8'b00000000;
		12'd1597: row_of_pixels <= 8'b00000000;
		12'd1598: row_of_pixels <= 8'b00000000;
		12'd1599: row_of_pixels <= 8'b00000000;
		12'd1600: row_of_pixels <= 8'b00000000;
		12'd1601: row_of_pixels <= 8'b00000000;
		12'd1602: row_of_pixels <= 8'b00111000;
		12'd1603: row_of_pixels <= 8'b00110000;
		12'd1604: row_of_pixels <= 8'b00110000;
		12'd1605: row_of_pixels <= 8'b00111100;
		12'd1606: row_of_pixels <= 8'b00110110;
		12'd1607: row_of_pixels <= 8'b00110011;
		12'd1608: row_of_pixels <= 8'b00110011;
		12'd1609: row_of_pixels <= 8'b00110011;
		12'd1610: row_of_pixels <= 8'b00110011;
		12'd1611: row_of_pixels <= 8'b01101110;
		12'd1612: row_of_pixels <= 8'b00000000;
		12'd1613: row_of_pixels <= 8'b00000000;
		12'd1614: row_of_pixels <= 8'b00000000;
		12'd1615: row_of_pixels <= 8'b00000000;
		12'd1616: row_of_pixels <= 8'b00000000;
		12'd1617: row_of_pixels <= 8'b00000000;
		12'd1618: row_of_pixels <= 8'b00000000;
		12'd1619: row_of_pixels <= 8'b00000000;
		12'd1620: row_of_pixels <= 8'b00000000;
		12'd1621: row_of_pixels <= 8'b00111110;
		12'd1622: row_of_pixels <= 8'b01100011;
		12'd1623: row_of_pixels <= 8'b01111111;
		12'd1624: row_of_pixels <= 8'b00000011;
		12'd1625: row_of_pixels <= 8'b00000011;
		12'd1626: row_of_pixels <= 8'b01100011;
		12'd1627: row_of_pixels <= 8'b00111110;
		12'd1628: row_of_pixels <= 8'b00000000;
		12'd1629: row_of_pixels <= 8'b00000000;
		12'd1630: row_of_pixels <= 8'b00000000;
		12'd1631: row_of_pixels <= 8'b00000000;
		12'd1632: row_of_pixels <= 8'b00000000;
		12'd1633: row_of_pixels <= 8'b00000000;
		12'd1634: row_of_pixels <= 8'b00011100;
		12'd1635: row_of_pixels <= 8'b00110110;
		12'd1636: row_of_pixels <= 8'b00100110;
		12'd1637: row_of_pixels <= 8'b00000110;
		12'd1638: row_of_pixels <= 8'b00001111;
		12'd1639: row_of_pixels <= 8'b00000110;
		12'd1640: row_of_pixels <= 8'b00000110;
		12'd1641: row_of_pixels <= 8'b00000110;
		12'd1642: row_of_pixels <= 8'b00000110;
		12'd1643: row_of_pixels <= 8'b00001111;
		12'd1644: row_of_pixels <= 8'b00000000;
		12'd1645: row_of_pixels <= 8'b00000000;
		12'd1646: row_of_pixels <= 8'b00000000;
		12'd1647: row_of_pixels <= 8'b00000000;
		12'd1648: row_of_pixels <= 8'b00000000;
		12'd1649: row_of_pixels <= 8'b00000000;
		12'd1650: row_of_pixels <= 8'b00000000;
		12'd1651: row_of_pixels <= 8'b00000000;
		12'd1652: row_of_pixels <= 8'b00000000;
		12'd1653: row_of_pixels <= 8'b01101110;
		12'd1654: row_of_pixels <= 8'b00110011;
		12'd1655: row_of_pixels <= 8'b00110011;
		12'd1656: row_of_pixels <= 8'b00110011;
		12'd1657: row_of_pixels <= 8'b00110011;
		12'd1658: row_of_pixels <= 8'b00110011;
		12'd1659: row_of_pixels <= 8'b00111110;
		12'd1660: row_of_pixels <= 8'b00110000;
		12'd1661: row_of_pixels <= 8'b00110011;
		12'd1662: row_of_pixels <= 8'b00011110;
		12'd1663: row_of_pixels <= 8'b00000000;
		12'd1664: row_of_pixels <= 8'b00000000;
		12'd1665: row_of_pixels <= 8'b00000000;
		12'd1666: row_of_pixels <= 8'b00000111;
		12'd1667: row_of_pixels <= 8'b00000110;
		12'd1668: row_of_pixels <= 8'b00000110;
		12'd1669: row_of_pixels <= 8'b00110110;
		12'd1670: row_of_pixels <= 8'b01101110;
		12'd1671: row_of_pixels <= 8'b01100110;
		12'd1672: row_of_pixels <= 8'b01100110;
		12'd1673: row_of_pixels <= 8'b01100110;
		12'd1674: row_of_pixels <= 8'b01100110;
		12'd1675: row_of_pixels <= 8'b01100111;
		12'd1676: row_of_pixels <= 8'b00000000;
		12'd1677: row_of_pixels <= 8'b00000000;
		12'd1678: row_of_pixels <= 8'b00000000;
		12'd1679: row_of_pixels <= 8'b00000000;
		12'd1680: row_of_pixels <= 8'b00000000;
		12'd1681: row_of_pixels <= 8'b00000000;
		12'd1682: row_of_pixels <= 8'b00011000;
		12'd1683: row_of_pixels <= 8'b00011000;
		12'd1684: row_of_pixels <= 8'b00000000;
		12'd1685: row_of_pixels <= 8'b00011100;
		12'd1686: row_of_pixels <= 8'b00011000;
		12'd1687: row_of_pixels <= 8'b00011000;
		12'd1688: row_of_pixels <= 8'b00011000;
		12'd1689: row_of_pixels <= 8'b00011000;
		12'd1690: row_of_pixels <= 8'b00011000;
		12'd1691: row_of_pixels <= 8'b00111100;
		12'd1692: row_of_pixels <= 8'b00000000;
		12'd1693: row_of_pixels <= 8'b00000000;
		12'd1694: row_of_pixels <= 8'b00000000;
		12'd1695: row_of_pixels <= 8'b00000000;
		12'd1696: row_of_pixels <= 8'b00000000;
		12'd1697: row_of_pixels <= 8'b00000000;
		12'd1698: row_of_pixels <= 8'b01100000;
		12'd1699: row_of_pixels <= 8'b01100000;
		12'd1700: row_of_pixels <= 8'b00000000;
		12'd1701: row_of_pixels <= 8'b01110000;
		12'd1702: row_of_pixels <= 8'b01100000;
		12'd1703: row_of_pixels <= 8'b01100000;
		12'd1704: row_of_pixels <= 8'b01100000;
		12'd1705: row_of_pixels <= 8'b01100000;
		12'd1706: row_of_pixels <= 8'b01100000;
		12'd1707: row_of_pixels <= 8'b01100000;
		12'd1708: row_of_pixels <= 8'b01100110;
		12'd1709: row_of_pixels <= 8'b01100110;
		12'd1710: row_of_pixels <= 8'b00111100;
		12'd1711: row_of_pixels <= 8'b00000000;
		12'd1712: row_of_pixels <= 8'b00000000;
		12'd1713: row_of_pixels <= 8'b00000000;
		12'd1714: row_of_pixels <= 8'b00000111;
		12'd1715: row_of_pixels <= 8'b00000110;
		12'd1716: row_of_pixels <= 8'b00000110;
		12'd1717: row_of_pixels <= 8'b01100110;
		12'd1718: row_of_pixels <= 8'b00110110;
		12'd1719: row_of_pixels <= 8'b00011110;
		12'd1720: row_of_pixels <= 8'b00011110;
		12'd1721: row_of_pixels <= 8'b00110110;
		12'd1722: row_of_pixels <= 8'b01100110;
		12'd1723: row_of_pixels <= 8'b01100111;
		12'd1724: row_of_pixels <= 8'b00000000;
		12'd1725: row_of_pixels <= 8'b00000000;
		12'd1726: row_of_pixels <= 8'b00000000;
		12'd1727: row_of_pixels <= 8'b00000000;
		12'd1728: row_of_pixels <= 8'b00000000;
		12'd1729: row_of_pixels <= 8'b00000000;
		12'd1730: row_of_pixels <= 8'b00011100;
		12'd1731: row_of_pixels <= 8'b00011000;
		12'd1732: row_of_pixels <= 8'b00011000;
		12'd1733: row_of_pixels <= 8'b00011000;
		12'd1734: row_of_pixels <= 8'b00011000;
		12'd1735: row_of_pixels <= 8'b00011000;
		12'd1736: row_of_pixels <= 8'b00011000;
		12'd1737: row_of_pixels <= 8'b00011000;
		12'd1738: row_of_pixels <= 8'b00011000;
		12'd1739: row_of_pixels <= 8'b00111100;
		12'd1740: row_of_pixels <= 8'b00000000;
		12'd1741: row_of_pixels <= 8'b00000000;
		12'd1742: row_of_pixels <= 8'b00000000;
		12'd1743: row_of_pixels <= 8'b00000000;
		12'd1744: row_of_pixels <= 8'b00000000;
		12'd1745: row_of_pixels <= 8'b00000000;
		12'd1746: row_of_pixels <= 8'b00000000;
		12'd1747: row_of_pixels <= 8'b00000000;
		12'd1748: row_of_pixels <= 8'b00000000;
		12'd1749: row_of_pixels <= 8'b01100111;
		12'd1750: row_of_pixels <= 8'b11111111;
		12'd1751: row_of_pixels <= 8'b11011011;
		12'd1752: row_of_pixels <= 8'b11011011;
		12'd1753: row_of_pixels <= 8'b11011011;
		12'd1754: row_of_pixels <= 8'b11011011;
		12'd1755: row_of_pixels <= 8'b11011011;
		12'd1756: row_of_pixels <= 8'b00000000;
		12'd1757: row_of_pixels <= 8'b00000000;
		12'd1758: row_of_pixels <= 8'b00000000;
		12'd1759: row_of_pixels <= 8'b00000000;
		12'd1760: row_of_pixels <= 8'b00000000;
		12'd1761: row_of_pixels <= 8'b00000000;
		12'd1762: row_of_pixels <= 8'b00000000;
		12'd1763: row_of_pixels <= 8'b00000000;
		12'd1764: row_of_pixels <= 8'b00000000;
		12'd1765: row_of_pixels <= 8'b00111011;
		12'd1766: row_of_pixels <= 8'b01100110;
		12'd1767: row_of_pixels <= 8'b01100110;
		12'd1768: row_of_pixels <= 8'b01100110;
		12'd1769: row_of_pixels <= 8'b01100110;
		12'd1770: row_of_pixels <= 8'b01100110;
		12'd1771: row_of_pixels <= 8'b01100110;
		12'd1772: row_of_pixels <= 8'b00000000;
		12'd1773: row_of_pixels <= 8'b00000000;
		12'd1774: row_of_pixels <= 8'b00000000;
		12'd1775: row_of_pixels <= 8'b00000000;
		12'd1776: row_of_pixels <= 8'b00000000;
		12'd1777: row_of_pixels <= 8'b00000000;
		12'd1778: row_of_pixels <= 8'b00000000;
		12'd1779: row_of_pixels <= 8'b00000000;
		12'd1780: row_of_pixels <= 8'b00000000;
		12'd1781: row_of_pixels <= 8'b00111110;
		12'd1782: row_of_pixels <= 8'b01100011;
		12'd1783: row_of_pixels <= 8'b01100011;
		12'd1784: row_of_pixels <= 8'b01100011;
		12'd1785: row_of_pixels <= 8'b01100011;
		12'd1786: row_of_pixels <= 8'b01100011;
		12'd1787: row_of_pixels <= 8'b00111110;
		12'd1788: row_of_pixels <= 8'b00000000;
		12'd1789: row_of_pixels <= 8'b00000000;
		12'd1790: row_of_pixels <= 8'b00000000;
		12'd1791: row_of_pixels <= 8'b00000000;
		12'd1792: row_of_pixels <= 8'b00000000;
		12'd1793: row_of_pixels <= 8'b00000000;
		12'd1794: row_of_pixels <= 8'b00000000;
		12'd1795: row_of_pixels <= 8'b00000000;
		12'd1796: row_of_pixels <= 8'b00000000;
		12'd1797: row_of_pixels <= 8'b00111011;
		12'd1798: row_of_pixels <= 8'b01100110;
		12'd1799: row_of_pixels <= 8'b01100110;
		12'd1800: row_of_pixels <= 8'b01100110;
		12'd1801: row_of_pixels <= 8'b01100110;
		12'd1802: row_of_pixels <= 8'b01100110;
		12'd1803: row_of_pixels <= 8'b00111110;
		12'd1804: row_of_pixels <= 8'b00000110;
		12'd1805: row_of_pixels <= 8'b00000110;
		12'd1806: row_of_pixels <= 8'b00001111;
		12'd1807: row_of_pixels <= 8'b00000000;
		12'd1808: row_of_pixels <= 8'b00000000;
		12'd1809: row_of_pixels <= 8'b00000000;
		12'd1810: row_of_pixels <= 8'b00000000;
		12'd1811: row_of_pixels <= 8'b00000000;
		12'd1812: row_of_pixels <= 8'b00000000;
		12'd1813: row_of_pixels <= 8'b01101110;
		12'd1814: row_of_pixels <= 8'b00110011;
		12'd1815: row_of_pixels <= 8'b00110011;
		12'd1816: row_of_pixels <= 8'b00110011;
		12'd1817: row_of_pixels <= 8'b00110011;
		12'd1818: row_of_pixels <= 8'b00110011;
		12'd1819: row_of_pixels <= 8'b00111110;
		12'd1820: row_of_pixels <= 8'b00110000;
		12'd1821: row_of_pixels <= 8'b00110000;
		12'd1822: row_of_pixels <= 8'b01111000;
		12'd1823: row_of_pixels <= 8'b00000000;
		12'd1824: row_of_pixels <= 8'b00000000;
		12'd1825: row_of_pixels <= 8'b00000000;
		12'd1826: row_of_pixels <= 8'b00000000;
		12'd1827: row_of_pixels <= 8'b00000000;
		12'd1828: row_of_pixels <= 8'b00000000;
		12'd1829: row_of_pixels <= 8'b00111011;
		12'd1830: row_of_pixels <= 8'b01101110;
		12'd1831: row_of_pixels <= 8'b01100110;
		12'd1832: row_of_pixels <= 8'b00000110;
		12'd1833: row_of_pixels <= 8'b00000110;
		12'd1834: row_of_pixels <= 8'b00000110;
		12'd1835: row_of_pixels <= 8'b00001111;
		12'd1836: row_of_pixels <= 8'b00000000;
		12'd1837: row_of_pixels <= 8'b00000000;
		12'd1838: row_of_pixels <= 8'b00000000;
		12'd1839: row_of_pixels <= 8'b00000000;
		12'd1840: row_of_pixels <= 8'b00000000;
		12'd1841: row_of_pixels <= 8'b00000000;
		12'd1842: row_of_pixels <= 8'b00000000;
		12'd1843: row_of_pixels <= 8'b00000000;
		12'd1844: row_of_pixels <= 8'b00000000;
		12'd1845: row_of_pixels <= 8'b00111110;
		12'd1846: row_of_pixels <= 8'b01100011;
		12'd1847: row_of_pixels <= 8'b00000110;
		12'd1848: row_of_pixels <= 8'b00011100;
		12'd1849: row_of_pixels <= 8'b00110000;
		12'd1850: row_of_pixels <= 8'b01100011;
		12'd1851: row_of_pixels <= 8'b00111110;
		12'd1852: row_of_pixels <= 8'b00000000;
		12'd1853: row_of_pixels <= 8'b00000000;
		12'd1854: row_of_pixels <= 8'b00000000;
		12'd1855: row_of_pixels <= 8'b00000000;
		12'd1856: row_of_pixels <= 8'b00000000;
		12'd1857: row_of_pixels <= 8'b00000000;
		12'd1858: row_of_pixels <= 8'b00001000;
		12'd1859: row_of_pixels <= 8'b00001100;
		12'd1860: row_of_pixels <= 8'b00001100;
		12'd1861: row_of_pixels <= 8'b00111111;
		12'd1862: row_of_pixels <= 8'b00001100;
		12'd1863: row_of_pixels <= 8'b00001100;
		12'd1864: row_of_pixels <= 8'b00001100;
		12'd1865: row_of_pixels <= 8'b00001100;
		12'd1866: row_of_pixels <= 8'b01101100;
		12'd1867: row_of_pixels <= 8'b00111000;
		12'd1868: row_of_pixels <= 8'b00000000;
		12'd1869: row_of_pixels <= 8'b00000000;
		12'd1870: row_of_pixels <= 8'b00000000;
		12'd1871: row_of_pixels <= 8'b00000000;
		12'd1872: row_of_pixels <= 8'b00000000;
		12'd1873: row_of_pixels <= 8'b00000000;
		12'd1874: row_of_pixels <= 8'b00000000;
		12'd1875: row_of_pixels <= 8'b00000000;
		12'd1876: row_of_pixels <= 8'b00000000;
		12'd1877: row_of_pixels <= 8'b00110011;
		12'd1878: row_of_pixels <= 8'b00110011;
		12'd1879: row_of_pixels <= 8'b00110011;
		12'd1880: row_of_pixels <= 8'b00110011;
		12'd1881: row_of_pixels <= 8'b00110011;
		12'd1882: row_of_pixels <= 8'b00110011;
		12'd1883: row_of_pixels <= 8'b01101110;
		12'd1884: row_of_pixels <= 8'b00000000;
		12'd1885: row_of_pixels <= 8'b00000000;
		12'd1886: row_of_pixels <= 8'b00000000;
		12'd1887: row_of_pixels <= 8'b00000000;
		12'd1888: row_of_pixels <= 8'b00000000;
		12'd1889: row_of_pixels <= 8'b00000000;
		12'd1890: row_of_pixels <= 8'b00000000;
		12'd1891: row_of_pixels <= 8'b00000000;
		12'd1892: row_of_pixels <= 8'b00000000;
		12'd1893: row_of_pixels <= 8'b11000011;
		12'd1894: row_of_pixels <= 8'b11000011;
		12'd1895: row_of_pixels <= 8'b11000011;
		12'd1896: row_of_pixels <= 8'b11000011;
		12'd1897: row_of_pixels <= 8'b01100110;
		12'd1898: row_of_pixels <= 8'b00111100;
		12'd1899: row_of_pixels <= 8'b00011000;
		12'd1900: row_of_pixels <= 8'b00000000;
		12'd1901: row_of_pixels <= 8'b00000000;
		12'd1902: row_of_pixels <= 8'b00000000;
		12'd1903: row_of_pixels <= 8'b00000000;
		12'd1904: row_of_pixels <= 8'b00000000;
		12'd1905: row_of_pixels <= 8'b00000000;
		12'd1906: row_of_pixels <= 8'b00000000;
		12'd1907: row_of_pixels <= 8'b00000000;
		12'd1908: row_of_pixels <= 8'b00000000;
		12'd1909: row_of_pixels <= 8'b11000011;
		12'd1910: row_of_pixels <= 8'b11000011;
		12'd1911: row_of_pixels <= 8'b11000011;
		12'd1912: row_of_pixels <= 8'b11011011;
		12'd1913: row_of_pixels <= 8'b11011011;
		12'd1914: row_of_pixels <= 8'b11111111;
		12'd1915: row_of_pixels <= 8'b01100110;
		12'd1916: row_of_pixels <= 8'b00000000;
		12'd1917: row_of_pixels <= 8'b00000000;
		12'd1918: row_of_pixels <= 8'b00000000;
		12'd1919: row_of_pixels <= 8'b00000000;
		12'd1920: row_of_pixels <= 8'b00000000;
		12'd1921: row_of_pixels <= 8'b00000000;
		12'd1922: row_of_pixels <= 8'b00000000;
		12'd1923: row_of_pixels <= 8'b00000000;
		12'd1924: row_of_pixels <= 8'b00000000;
		12'd1925: row_of_pixels <= 8'b11000011;
		12'd1926: row_of_pixels <= 8'b01100110;
		12'd1927: row_of_pixels <= 8'b00111100;
		12'd1928: row_of_pixels <= 8'b00011000;
		12'd1929: row_of_pixels <= 8'b00111100;
		12'd1930: row_of_pixels <= 8'b01100110;
		12'd1931: row_of_pixels <= 8'b11000011;
		12'd1932: row_of_pixels <= 8'b00000000;
		12'd1933: row_of_pixels <= 8'b00000000;
		12'd1934: row_of_pixels <= 8'b00000000;
		12'd1935: row_of_pixels <= 8'b00000000;
		12'd1936: row_of_pixels <= 8'b00000000;
		12'd1937: row_of_pixels <= 8'b00000000;
		12'd1938: row_of_pixels <= 8'b00000000;
		12'd1939: row_of_pixels <= 8'b00000000;
		12'd1940: row_of_pixels <= 8'b00000000;
		12'd1941: row_of_pixels <= 8'b01100011;
		12'd1942: row_of_pixels <= 8'b01100011;
		12'd1943: row_of_pixels <= 8'b01100011;
		12'd1944: row_of_pixels <= 8'b01100011;
		12'd1945: row_of_pixels <= 8'b01100011;
		12'd1946: row_of_pixels <= 8'b01100011;
		12'd1947: row_of_pixels <= 8'b01111110;
		12'd1948: row_of_pixels <= 8'b01100000;
		12'd1949: row_of_pixels <= 8'b00110000;
		12'd1950: row_of_pixels <= 8'b00011111;
		12'd1951: row_of_pixels <= 8'b00000000;
		12'd1952: row_of_pixels <= 8'b00000000;
		12'd1953: row_of_pixels <= 8'b00000000;
		12'd1954: row_of_pixels <= 8'b00000000;
		12'd1955: row_of_pixels <= 8'b00000000;
		12'd1956: row_of_pixels <= 8'b00000000;
		12'd1957: row_of_pixels <= 8'b01111111;
		12'd1958: row_of_pixels <= 8'b00110011;
		12'd1959: row_of_pixels <= 8'b00011000;
		12'd1960: row_of_pixels <= 8'b00001100;
		12'd1961: row_of_pixels <= 8'b00000110;
		12'd1962: row_of_pixels <= 8'b01100011;
		12'd1963: row_of_pixels <= 8'b01111111;
		12'd1964: row_of_pixels <= 8'b00000000;
		12'd1965: row_of_pixels <= 8'b00000000;
		12'd1966: row_of_pixels <= 8'b00000000;
		12'd1967: row_of_pixels <= 8'b00000000;
		12'd1968: row_of_pixels <= 8'b00000000;
		12'd1969: row_of_pixels <= 8'b00000000;
		12'd1970: row_of_pixels <= 8'b01110000;
		12'd1971: row_of_pixels <= 8'b00011000;
		12'd1972: row_of_pixels <= 8'b00011000;
		12'd1973: row_of_pixels <= 8'b00011000;
		12'd1974: row_of_pixels <= 8'b00001110;
		12'd1975: row_of_pixels <= 8'b00011000;
		12'd1976: row_of_pixels <= 8'b00011000;
		12'd1977: row_of_pixels <= 8'b00011000;
		12'd1978: row_of_pixels <= 8'b00011000;
		12'd1979: row_of_pixels <= 8'b01110000;
		12'd1980: row_of_pixels <= 8'b00000000;
		12'd1981: row_of_pixels <= 8'b00000000;
		12'd1982: row_of_pixels <= 8'b00000000;
		12'd1983: row_of_pixels <= 8'b00000000;
		12'd1984: row_of_pixels <= 8'b00000000;
		12'd1985: row_of_pixels <= 8'b00000000;
		12'd1986: row_of_pixels <= 8'b00011000;
		12'd1987: row_of_pixels <= 8'b00011000;
		12'd1988: row_of_pixels <= 8'b00011000;
		12'd1989: row_of_pixels <= 8'b00011000;
		12'd1990: row_of_pixels <= 8'b00000000;
		12'd1991: row_of_pixels <= 8'b00011000;
		12'd1992: row_of_pixels <= 8'b00011000;
		12'd1993: row_of_pixels <= 8'b00011000;
		12'd1994: row_of_pixels <= 8'b00011000;
		12'd1995: row_of_pixels <= 8'b00011000;
		12'd1996: row_of_pixels <= 8'b00000000;
		12'd1997: row_of_pixels <= 8'b00000000;
		12'd1998: row_of_pixels <= 8'b00000000;
		12'd1999: row_of_pixels <= 8'b00000000;
		12'd2000: row_of_pixels <= 8'b00000000;
		12'd2001: row_of_pixels <= 8'b00000000;
		12'd2002: row_of_pixels <= 8'b00001110;
		12'd2003: row_of_pixels <= 8'b00011000;
		12'd2004: row_of_pixels <= 8'b00011000;
		12'd2005: row_of_pixels <= 8'b00011000;
		12'd2006: row_of_pixels <= 8'b01110000;
		12'd2007: row_of_pixels <= 8'b00011000;
		12'd2008: row_of_pixels <= 8'b00011000;
		12'd2009: row_of_pixels <= 8'b00011000;
		12'd2010: row_of_pixels <= 8'b00011000;
		12'd2011: row_of_pixels <= 8'b00001110;
		12'd2012: row_of_pixels <= 8'b00000000;
		12'd2013: row_of_pixels <= 8'b00000000;
		12'd2014: row_of_pixels <= 8'b00000000;
		12'd2015: row_of_pixels <= 8'b00000000;
		12'd2016: row_of_pixels <= 8'b00000000;
		12'd2017: row_of_pixels <= 8'b00000000;
		12'd2018: row_of_pixels <= 8'b01101110;
		12'd2019: row_of_pixels <= 8'b00111011;
		12'd2020: row_of_pixels <= 8'b00000000;
		12'd2021: row_of_pixels <= 8'b00000000;
		12'd2022: row_of_pixels <= 8'b00000000;
		12'd2023: row_of_pixels <= 8'b00000000;
		12'd2024: row_of_pixels <= 8'b00000000;
		12'd2025: row_of_pixels <= 8'b00000000;
		12'd2026: row_of_pixels <= 8'b00000000;
		12'd2027: row_of_pixels <= 8'b00000000;
		12'd2028: row_of_pixels <= 8'b00000000;
		12'd2029: row_of_pixels <= 8'b00000000;
		12'd2030: row_of_pixels <= 8'b00000000;
		12'd2031: row_of_pixels <= 8'b00000000;
		12'd2032: row_of_pixels <= 8'b00000000;
		12'd2033: row_of_pixels <= 8'b00000000;
		12'd2034: row_of_pixels <= 8'b00000000;
		12'd2035: row_of_pixels <= 8'b00000000;
		12'd2036: row_of_pixels <= 8'b00001000;
		12'd2037: row_of_pixels <= 8'b00011100;
		12'd2038: row_of_pixels <= 8'b00110110;
		12'd2039: row_of_pixels <= 8'b01100011;
		12'd2040: row_of_pixels <= 8'b01100011;
		12'd2041: row_of_pixels <= 8'b01100011;
		12'd2042: row_of_pixels <= 8'b01111111;
		12'd2043: row_of_pixels <= 8'b00000000;
		12'd2044: row_of_pixels <= 8'b00000000;
		12'd2045: row_of_pixels <= 8'b00000000;
		12'd2046: row_of_pixels <= 8'b00000000;
		12'd2047: row_of_pixels <= 8'b00000000;
		12'd2048: row_of_pixels <= 8'b00000000;
		12'd2049: row_of_pixels <= 8'b00000000;
		12'd2050: row_of_pixels <= 8'b00111100;
		12'd2051: row_of_pixels <= 8'b01100110;
		12'd2052: row_of_pixels <= 8'b01000011;
		12'd2053: row_of_pixels <= 8'b00000011;
		12'd2054: row_of_pixels <= 8'b00000011;
		12'd2055: row_of_pixels <= 8'b00000011;
		12'd2056: row_of_pixels <= 8'b01000011;
		12'd2057: row_of_pixels <= 8'b01100110;
		12'd2058: row_of_pixels <= 8'b00111100;
		12'd2059: row_of_pixels <= 8'b00110000;
		12'd2060: row_of_pixels <= 8'b01100000;
		12'd2061: row_of_pixels <= 8'b00111110;
		12'd2062: row_of_pixels <= 8'b00000000;
		12'd2063: row_of_pixels <= 8'b00000000;
		12'd2064: row_of_pixels <= 8'b00000000;
		12'd2065: row_of_pixels <= 8'b00000000;
		12'd2066: row_of_pixels <= 8'b00110011;
		12'd2067: row_of_pixels <= 8'b00000000;
		12'd2068: row_of_pixels <= 8'b00000000;
		12'd2069: row_of_pixels <= 8'b00110011;
		12'd2070: row_of_pixels <= 8'b00110011;
		12'd2071: row_of_pixels <= 8'b00110011;
		12'd2072: row_of_pixels <= 8'b00110011;
		12'd2073: row_of_pixels <= 8'b00110011;
		12'd2074: row_of_pixels <= 8'b00110011;
		12'd2075: row_of_pixels <= 8'b01101110;
		12'd2076: row_of_pixels <= 8'b00000000;
		12'd2077: row_of_pixels <= 8'b00000000;
		12'd2078: row_of_pixels <= 8'b00000000;
		12'd2079: row_of_pixels <= 8'b00000000;
		12'd2080: row_of_pixels <= 8'b00000000;
		12'd2081: row_of_pixels <= 8'b00110000;
		12'd2082: row_of_pixels <= 8'b00011000;
		12'd2083: row_of_pixels <= 8'b00001100;
		12'd2084: row_of_pixels <= 8'b00000000;
		12'd2085: row_of_pixels <= 8'b00111110;
		12'd2086: row_of_pixels <= 8'b01100011;
		12'd2087: row_of_pixels <= 8'b01111111;
		12'd2088: row_of_pixels <= 8'b00000011;
		12'd2089: row_of_pixels <= 8'b00000011;
		12'd2090: row_of_pixels <= 8'b01100011;
		12'd2091: row_of_pixels <= 8'b00111110;
		12'd2092: row_of_pixels <= 8'b00000000;
		12'd2093: row_of_pixels <= 8'b00000000;
		12'd2094: row_of_pixels <= 8'b00000000;
		12'd2095: row_of_pixels <= 8'b00000000;
		12'd2096: row_of_pixels <= 8'b00000000;
		12'd2097: row_of_pixels <= 8'b00001000;
		12'd2098: row_of_pixels <= 8'b00011100;
		12'd2099: row_of_pixels <= 8'b00110110;
		12'd2100: row_of_pixels <= 8'b00000000;
		12'd2101: row_of_pixels <= 8'b00011110;
		12'd2102: row_of_pixels <= 8'b00110000;
		12'd2103: row_of_pixels <= 8'b00111110;
		12'd2104: row_of_pixels <= 8'b00110011;
		12'd2105: row_of_pixels <= 8'b00110011;
		12'd2106: row_of_pixels <= 8'b00110011;
		12'd2107: row_of_pixels <= 8'b01101110;
		12'd2108: row_of_pixels <= 8'b00000000;
		12'd2109: row_of_pixels <= 8'b00000000;
		12'd2110: row_of_pixels <= 8'b00000000;
		12'd2111: row_of_pixels <= 8'b00000000;
		12'd2112: row_of_pixels <= 8'b00000000;
		12'd2113: row_of_pixels <= 8'b00000000;
		12'd2114: row_of_pixels <= 8'b00110011;
		12'd2115: row_of_pixels <= 8'b00000000;
		12'd2116: row_of_pixels <= 8'b00000000;
		12'd2117: row_of_pixels <= 8'b00011110;
		12'd2118: row_of_pixels <= 8'b00110000;
		12'd2119: row_of_pixels <= 8'b00111110;
		12'd2120: row_of_pixels <= 8'b00110011;
		12'd2121: row_of_pixels <= 8'b00110011;
		12'd2122: row_of_pixels <= 8'b00110011;
		12'd2123: row_of_pixels <= 8'b01101110;
		12'd2124: row_of_pixels <= 8'b00000000;
		12'd2125: row_of_pixels <= 8'b00000000;
		12'd2126: row_of_pixels <= 8'b00000000;
		12'd2127: row_of_pixels <= 8'b00000000;
		12'd2128: row_of_pixels <= 8'b00000000;
		12'd2129: row_of_pixels <= 8'b00000110;
		12'd2130: row_of_pixels <= 8'b00001100;
		12'd2131: row_of_pixels <= 8'b00011000;
		12'd2132: row_of_pixels <= 8'b00000000;
		12'd2133: row_of_pixels <= 8'b00011110;
		12'd2134: row_of_pixels <= 8'b00110000;
		12'd2135: row_of_pixels <= 8'b00111110;
		12'd2136: row_of_pixels <= 8'b00110011;
		12'd2137: row_of_pixels <= 8'b00110011;
		12'd2138: row_of_pixels <= 8'b00110011;
		12'd2139: row_of_pixels <= 8'b01101110;
		12'd2140: row_of_pixels <= 8'b00000000;
		12'd2141: row_of_pixels <= 8'b00000000;
		12'd2142: row_of_pixels <= 8'b00000000;
		12'd2143: row_of_pixels <= 8'b00000000;
		12'd2144: row_of_pixels <= 8'b00000000;
		12'd2145: row_of_pixels <= 8'b00011100;
		12'd2146: row_of_pixels <= 8'b00110110;
		12'd2147: row_of_pixels <= 8'b00011100;
		12'd2148: row_of_pixels <= 8'b00000000;
		12'd2149: row_of_pixels <= 8'b00011110;
		12'd2150: row_of_pixels <= 8'b00110000;
		12'd2151: row_of_pixels <= 8'b00111110;
		12'd2152: row_of_pixels <= 8'b00110011;
		12'd2153: row_of_pixels <= 8'b00110011;
		12'd2154: row_of_pixels <= 8'b00110011;
		12'd2155: row_of_pixels <= 8'b01101110;
		12'd2156: row_of_pixels <= 8'b00000000;
		12'd2157: row_of_pixels <= 8'b00000000;
		12'd2158: row_of_pixels <= 8'b00000000;
		12'd2159: row_of_pixels <= 8'b00000000;
		12'd2160: row_of_pixels <= 8'b00000000;
		12'd2161: row_of_pixels <= 8'b00000000;
		12'd2162: row_of_pixels <= 8'b00000000;
		12'd2163: row_of_pixels <= 8'b00000000;
		12'd2164: row_of_pixels <= 8'b00111100;
		12'd2165: row_of_pixels <= 8'b01100110;
		12'd2166: row_of_pixels <= 8'b00000110;
		12'd2167: row_of_pixels <= 8'b00000110;
		12'd2168: row_of_pixels <= 8'b01100110;
		12'd2169: row_of_pixels <= 8'b00111100;
		12'd2170: row_of_pixels <= 8'b00110000;
		12'd2171: row_of_pixels <= 8'b01100000;
		12'd2172: row_of_pixels <= 8'b00111100;
		12'd2173: row_of_pixels <= 8'b00000000;
		12'd2174: row_of_pixels <= 8'b00000000;
		12'd2175: row_of_pixels <= 8'b00000000;
		12'd2176: row_of_pixels <= 8'b00000000;
		12'd2177: row_of_pixels <= 8'b00001000;
		12'd2178: row_of_pixels <= 8'b00011100;
		12'd2179: row_of_pixels <= 8'b00110110;
		12'd2180: row_of_pixels <= 8'b00000000;
		12'd2181: row_of_pixels <= 8'b00111110;
		12'd2182: row_of_pixels <= 8'b01100011;
		12'd2183: row_of_pixels <= 8'b01111111;
		12'd2184: row_of_pixels <= 8'b00000011;
		12'd2185: row_of_pixels <= 8'b00000011;
		12'd2186: row_of_pixels <= 8'b01100011;
		12'd2187: row_of_pixels <= 8'b00111110;
		12'd2188: row_of_pixels <= 8'b00000000;
		12'd2189: row_of_pixels <= 8'b00000000;
		12'd2190: row_of_pixels <= 8'b00000000;
		12'd2191: row_of_pixels <= 8'b00000000;
		12'd2192: row_of_pixels <= 8'b00000000;
		12'd2193: row_of_pixels <= 8'b00000000;
		12'd2194: row_of_pixels <= 8'b01100011;
		12'd2195: row_of_pixels <= 8'b00000000;
		12'd2196: row_of_pixels <= 8'b00000000;
		12'd2197: row_of_pixels <= 8'b00111110;
		12'd2198: row_of_pixels <= 8'b01100011;
		12'd2199: row_of_pixels <= 8'b01111111;
		12'd2200: row_of_pixels <= 8'b00000011;
		12'd2201: row_of_pixels <= 8'b00000011;
		12'd2202: row_of_pixels <= 8'b01100011;
		12'd2203: row_of_pixels <= 8'b00111110;
		12'd2204: row_of_pixels <= 8'b00000000;
		12'd2205: row_of_pixels <= 8'b00000000;
		12'd2206: row_of_pixels <= 8'b00000000;
		12'd2207: row_of_pixels <= 8'b00000000;
		12'd2208: row_of_pixels <= 8'b00000000;
		12'd2209: row_of_pixels <= 8'b00000110;
		12'd2210: row_of_pixels <= 8'b00001100;
		12'd2211: row_of_pixels <= 8'b00011000;
		12'd2212: row_of_pixels <= 8'b00000000;
		12'd2213: row_of_pixels <= 8'b00111110;
		12'd2214: row_of_pixels <= 8'b01100011;
		12'd2215: row_of_pixels <= 8'b01111111;
		12'd2216: row_of_pixels <= 8'b00000011;
		12'd2217: row_of_pixels <= 8'b00000011;
		12'd2218: row_of_pixels <= 8'b01100011;
		12'd2219: row_of_pixels <= 8'b00111110;
		12'd2220: row_of_pixels <= 8'b00000000;
		12'd2221: row_of_pixels <= 8'b00000000;
		12'd2222: row_of_pixels <= 8'b00000000;
		12'd2223: row_of_pixels <= 8'b00000000;
		12'd2224: row_of_pixels <= 8'b00000000;
		12'd2225: row_of_pixels <= 8'b00000000;
		12'd2226: row_of_pixels <= 8'b01100110;
		12'd2227: row_of_pixels <= 8'b00000000;
		12'd2228: row_of_pixels <= 8'b00000000;
		12'd2229: row_of_pixels <= 8'b00011100;
		12'd2230: row_of_pixels <= 8'b00011000;
		12'd2231: row_of_pixels <= 8'b00011000;
		12'd2232: row_of_pixels <= 8'b00011000;
		12'd2233: row_of_pixels <= 8'b00011000;
		12'd2234: row_of_pixels <= 8'b00011000;
		12'd2235: row_of_pixels <= 8'b00111100;
		12'd2236: row_of_pixels <= 8'b00000000;
		12'd2237: row_of_pixels <= 8'b00000000;
		12'd2238: row_of_pixels <= 8'b00000000;
		12'd2239: row_of_pixels <= 8'b00000000;
		12'd2240: row_of_pixels <= 8'b00000000;
		12'd2241: row_of_pixels <= 8'b00011000;
		12'd2242: row_of_pixels <= 8'b00111100;
		12'd2243: row_of_pixels <= 8'b01100110;
		12'd2244: row_of_pixels <= 8'b00000000;
		12'd2245: row_of_pixels <= 8'b00011100;
		12'd2246: row_of_pixels <= 8'b00011000;
		12'd2247: row_of_pixels <= 8'b00011000;
		12'd2248: row_of_pixels <= 8'b00011000;
		12'd2249: row_of_pixels <= 8'b00011000;
		12'd2250: row_of_pixels <= 8'b00011000;
		12'd2251: row_of_pixels <= 8'b00111100;
		12'd2252: row_of_pixels <= 8'b00000000;
		12'd2253: row_of_pixels <= 8'b00000000;
		12'd2254: row_of_pixels <= 8'b00000000;
		12'd2255: row_of_pixels <= 8'b00000000;
		12'd2256: row_of_pixels <= 8'b00000000;
		12'd2257: row_of_pixels <= 8'b00000110;
		12'd2258: row_of_pixels <= 8'b00001100;
		12'd2259: row_of_pixels <= 8'b00011000;
		12'd2260: row_of_pixels <= 8'b00000000;
		12'd2261: row_of_pixels <= 8'b00011100;
		12'd2262: row_of_pixels <= 8'b00011000;
		12'd2263: row_of_pixels <= 8'b00011000;
		12'd2264: row_of_pixels <= 8'b00011000;
		12'd2265: row_of_pixels <= 8'b00011000;
		12'd2266: row_of_pixels <= 8'b00011000;
		12'd2267: row_of_pixels <= 8'b00111100;
		12'd2268: row_of_pixels <= 8'b00000000;
		12'd2269: row_of_pixels <= 8'b00000000;
		12'd2270: row_of_pixels <= 8'b00000000;
		12'd2271: row_of_pixels <= 8'b00000000;
		12'd2272: row_of_pixels <= 8'b00000000;
		12'd2273: row_of_pixels <= 8'b01100011;
		12'd2274: row_of_pixels <= 8'b00000000;
		12'd2275: row_of_pixels <= 8'b00001000;
		12'd2276: row_of_pixels <= 8'b00011100;
		12'd2277: row_of_pixels <= 8'b00110110;
		12'd2278: row_of_pixels <= 8'b01100011;
		12'd2279: row_of_pixels <= 8'b01100011;
		12'd2280: row_of_pixels <= 8'b01111111;
		12'd2281: row_of_pixels <= 8'b01100011;
		12'd2282: row_of_pixels <= 8'b01100011;
		12'd2283: row_of_pixels <= 8'b01100011;
		12'd2284: row_of_pixels <= 8'b00000000;
		12'd2285: row_of_pixels <= 8'b00000000;
		12'd2286: row_of_pixels <= 8'b00000000;
		12'd2287: row_of_pixels <= 8'b00000000;
		12'd2288: row_of_pixels <= 8'b00011100;
		12'd2289: row_of_pixels <= 8'b00110110;
		12'd2290: row_of_pixels <= 8'b00011100;
		12'd2291: row_of_pixels <= 8'b00000000;
		12'd2292: row_of_pixels <= 8'b00011100;
		12'd2293: row_of_pixels <= 8'b00110110;
		12'd2294: row_of_pixels <= 8'b01100011;
		12'd2295: row_of_pixels <= 8'b01100011;
		12'd2296: row_of_pixels <= 8'b01111111;
		12'd2297: row_of_pixels <= 8'b01100011;
		12'd2298: row_of_pixels <= 8'b01100011;
		12'd2299: row_of_pixels <= 8'b01100011;
		12'd2300: row_of_pixels <= 8'b00000000;
		12'd2301: row_of_pixels <= 8'b00000000;
		12'd2302: row_of_pixels <= 8'b00000000;
		12'd2303: row_of_pixels <= 8'b00000000;
		12'd2304: row_of_pixels <= 8'b00011000;
		12'd2305: row_of_pixels <= 8'b00001100;
		12'd2306: row_of_pixels <= 8'b00000110;
		12'd2307: row_of_pixels <= 8'b00000000;
		12'd2308: row_of_pixels <= 8'b01111111;
		12'd2309: row_of_pixels <= 8'b01100110;
		12'd2310: row_of_pixels <= 8'b00000110;
		12'd2311: row_of_pixels <= 8'b00111110;
		12'd2312: row_of_pixels <= 8'b00000110;
		12'd2313: row_of_pixels <= 8'b00000110;
		12'd2314: row_of_pixels <= 8'b01100110;
		12'd2315: row_of_pixels <= 8'b01111111;
		12'd2316: row_of_pixels <= 8'b00000000;
		12'd2317: row_of_pixels <= 8'b00000000;
		12'd2318: row_of_pixels <= 8'b00000000;
		12'd2319: row_of_pixels <= 8'b00000000;
		12'd2320: row_of_pixels <= 8'b00000000;
		12'd2321: row_of_pixels <= 8'b00000000;
		12'd2322: row_of_pixels <= 8'b00000000;
		12'd2323: row_of_pixels <= 8'b00000000;
		12'd2324: row_of_pixels <= 8'b00000000;
		12'd2325: row_of_pixels <= 8'b01110110;
		12'd2326: row_of_pixels <= 8'b11011100;
		12'd2327: row_of_pixels <= 8'b11011000;
		12'd2328: row_of_pixels <= 8'b01111110;
		12'd2329: row_of_pixels <= 8'b00011011;
		12'd2330: row_of_pixels <= 8'b00111011;
		12'd2331: row_of_pixels <= 8'b11101110;
		12'd2332: row_of_pixels <= 8'b00000000;
		12'd2333: row_of_pixels <= 8'b00000000;
		12'd2334: row_of_pixels <= 8'b00000000;
		12'd2335: row_of_pixels <= 8'b00000000;
		12'd2336: row_of_pixels <= 8'b00000000;
		12'd2337: row_of_pixels <= 8'b00000000;
		12'd2338: row_of_pixels <= 8'b01111100;
		12'd2339: row_of_pixels <= 8'b00110110;
		12'd2340: row_of_pixels <= 8'b00110011;
		12'd2341: row_of_pixels <= 8'b00110011;
		12'd2342: row_of_pixels <= 8'b01111111;
		12'd2343: row_of_pixels <= 8'b00110011;
		12'd2344: row_of_pixels <= 8'b00110011;
		12'd2345: row_of_pixels <= 8'b00110011;
		12'd2346: row_of_pixels <= 8'b00110011;
		12'd2347: row_of_pixels <= 8'b01110011;
		12'd2348: row_of_pixels <= 8'b00000000;
		12'd2349: row_of_pixels <= 8'b00000000;
		12'd2350: row_of_pixels <= 8'b00000000;
		12'd2351: row_of_pixels <= 8'b00000000;
		12'd2352: row_of_pixels <= 8'b00000000;
		12'd2353: row_of_pixels <= 8'b00001000;
		12'd2354: row_of_pixels <= 8'b00011100;
		12'd2355: row_of_pixels <= 8'b00110110;
		12'd2356: row_of_pixels <= 8'b00000000;
		12'd2357: row_of_pixels <= 8'b00111110;
		12'd2358: row_of_pixels <= 8'b01100011;
		12'd2359: row_of_pixels <= 8'b01100011;
		12'd2360: row_of_pixels <= 8'b01100011;
		12'd2361: row_of_pixels <= 8'b01100011;
		12'd2362: row_of_pixels <= 8'b01100011;
		12'd2363: row_of_pixels <= 8'b00111110;
		12'd2364: row_of_pixels <= 8'b00000000;
		12'd2365: row_of_pixels <= 8'b00000000;
		12'd2366: row_of_pixels <= 8'b00000000;
		12'd2367: row_of_pixels <= 8'b00000000;
		12'd2368: row_of_pixels <= 8'b00000000;
		12'd2369: row_of_pixels <= 8'b00000000;
		12'd2370: row_of_pixels <= 8'b01100011;
		12'd2371: row_of_pixels <= 8'b00000000;
		12'd2372: row_of_pixels <= 8'b00000000;
		12'd2373: row_of_pixels <= 8'b00111110;
		12'd2374: row_of_pixels <= 8'b01100011;
		12'd2375: row_of_pixels <= 8'b01100011;
		12'd2376: row_of_pixels <= 8'b01100011;
		12'd2377: row_of_pixels <= 8'b01100011;
		12'd2378: row_of_pixels <= 8'b01100011;
		12'd2379: row_of_pixels <= 8'b00111110;
		12'd2380: row_of_pixels <= 8'b00000000;
		12'd2381: row_of_pixels <= 8'b00000000;
		12'd2382: row_of_pixels <= 8'b00000000;
		12'd2383: row_of_pixels <= 8'b00000000;
		12'd2384: row_of_pixels <= 8'b00000000;
		12'd2385: row_of_pixels <= 8'b00000110;
		12'd2386: row_of_pixels <= 8'b00001100;
		12'd2387: row_of_pixels <= 8'b00011000;
		12'd2388: row_of_pixels <= 8'b00000000;
		12'd2389: row_of_pixels <= 8'b00111110;
		12'd2390: row_of_pixels <= 8'b01100011;
		12'd2391: row_of_pixels <= 8'b01100011;
		12'd2392: row_of_pixels <= 8'b01100011;
		12'd2393: row_of_pixels <= 8'b01100011;
		12'd2394: row_of_pixels <= 8'b01100011;
		12'd2395: row_of_pixels <= 8'b00111110;
		12'd2396: row_of_pixels <= 8'b00000000;
		12'd2397: row_of_pixels <= 8'b00000000;
		12'd2398: row_of_pixels <= 8'b00000000;
		12'd2399: row_of_pixels <= 8'b00000000;
		12'd2400: row_of_pixels <= 8'b00000000;
		12'd2401: row_of_pixels <= 8'b00001100;
		12'd2402: row_of_pixels <= 8'b00011110;
		12'd2403: row_of_pixels <= 8'b00110011;
		12'd2404: row_of_pixels <= 8'b00000000;
		12'd2405: row_of_pixels <= 8'b00110011;
		12'd2406: row_of_pixels <= 8'b00110011;
		12'd2407: row_of_pixels <= 8'b00110011;
		12'd2408: row_of_pixels <= 8'b00110011;
		12'd2409: row_of_pixels <= 8'b00110011;
		12'd2410: row_of_pixels <= 8'b00110011;
		12'd2411: row_of_pixels <= 8'b01101110;
		12'd2412: row_of_pixels <= 8'b00000000;
		12'd2413: row_of_pixels <= 8'b00000000;
		12'd2414: row_of_pixels <= 8'b00000000;
		12'd2415: row_of_pixels <= 8'b00000000;
		12'd2416: row_of_pixels <= 8'b00000000;
		12'd2417: row_of_pixels <= 8'b00000110;
		12'd2418: row_of_pixels <= 8'b00001100;
		12'd2419: row_of_pixels <= 8'b00011000;
		12'd2420: row_of_pixels <= 8'b00000000;
		12'd2421: row_of_pixels <= 8'b00110011;
		12'd2422: row_of_pixels <= 8'b00110011;
		12'd2423: row_of_pixels <= 8'b00110011;
		12'd2424: row_of_pixels <= 8'b00110011;
		12'd2425: row_of_pixels <= 8'b00110011;
		12'd2426: row_of_pixels <= 8'b00110011;
		12'd2427: row_of_pixels <= 8'b01101110;
		12'd2428: row_of_pixels <= 8'b00000000;
		12'd2429: row_of_pixels <= 8'b00000000;
		12'd2430: row_of_pixels <= 8'b00000000;
		12'd2431: row_of_pixels <= 8'b00000000;
		12'd2432: row_of_pixels <= 8'b00000000;
		12'd2433: row_of_pixels <= 8'b00000000;
		12'd2434: row_of_pixels <= 8'b01100011;
		12'd2435: row_of_pixels <= 8'b00000000;
		12'd2436: row_of_pixels <= 8'b00000000;
		12'd2437: row_of_pixels <= 8'b01100011;
		12'd2438: row_of_pixels <= 8'b01100011;
		12'd2439: row_of_pixels <= 8'b01100011;
		12'd2440: row_of_pixels <= 8'b01100011;
		12'd2441: row_of_pixels <= 8'b01100011;
		12'd2442: row_of_pixels <= 8'b01100011;
		12'd2443: row_of_pixels <= 8'b01111110;
		12'd2444: row_of_pixels <= 8'b01100000;
		12'd2445: row_of_pixels <= 8'b00110000;
		12'd2446: row_of_pixels <= 8'b00011110;
		12'd2447: row_of_pixels <= 8'b00000000;
		12'd2448: row_of_pixels <= 8'b00000000;
		12'd2449: row_of_pixels <= 8'b01100011;
		12'd2450: row_of_pixels <= 8'b00000000;
		12'd2451: row_of_pixels <= 8'b00111110;
		12'd2452: row_of_pixels <= 8'b01100011;
		12'd2453: row_of_pixels <= 8'b01100011;
		12'd2454: row_of_pixels <= 8'b01100011;
		12'd2455: row_of_pixels <= 8'b01100011;
		12'd2456: row_of_pixels <= 8'b01100011;
		12'd2457: row_of_pixels <= 8'b01100011;
		12'd2458: row_of_pixels <= 8'b01100011;
		12'd2459: row_of_pixels <= 8'b00111110;
		12'd2460: row_of_pixels <= 8'b00000000;
		12'd2461: row_of_pixels <= 8'b00000000;
		12'd2462: row_of_pixels <= 8'b00000000;
		12'd2463: row_of_pixels <= 8'b00000000;
		12'd2464: row_of_pixels <= 8'b00000000;
		12'd2465: row_of_pixels <= 8'b01100011;
		12'd2466: row_of_pixels <= 8'b00000000;
		12'd2467: row_of_pixels <= 8'b01100011;
		12'd2468: row_of_pixels <= 8'b01100011;
		12'd2469: row_of_pixels <= 8'b01100011;
		12'd2470: row_of_pixels <= 8'b01100011;
		12'd2471: row_of_pixels <= 8'b01100011;
		12'd2472: row_of_pixels <= 8'b01100011;
		12'd2473: row_of_pixels <= 8'b01100011;
		12'd2474: row_of_pixels <= 8'b01100011;
		12'd2475: row_of_pixels <= 8'b00111110;
		12'd2476: row_of_pixels <= 8'b00000000;
		12'd2477: row_of_pixels <= 8'b00000000;
		12'd2478: row_of_pixels <= 8'b00000000;
		12'd2479: row_of_pixels <= 8'b00000000;
		12'd2480: row_of_pixels <= 8'b00000000;
		12'd2481: row_of_pixels <= 8'b00011000;
		12'd2482: row_of_pixels <= 8'b00011000;
		12'd2483: row_of_pixels <= 8'b01111110;
		12'd2484: row_of_pixels <= 8'b11000011;
		12'd2485: row_of_pixels <= 8'b00000011;
		12'd2486: row_of_pixels <= 8'b00000011;
		12'd2487: row_of_pixels <= 8'b00000011;
		12'd2488: row_of_pixels <= 8'b11000011;
		12'd2489: row_of_pixels <= 8'b01111110;
		12'd2490: row_of_pixels <= 8'b00011000;
		12'd2491: row_of_pixels <= 8'b00011000;
		12'd2492: row_of_pixels <= 8'b00000000;
		12'd2493: row_of_pixels <= 8'b00000000;
		12'd2494: row_of_pixels <= 8'b00000000;
		12'd2495: row_of_pixels <= 8'b00000000;
		12'd2496: row_of_pixels <= 8'b00000000;
		12'd2497: row_of_pixels <= 8'b00011100;
		12'd2498: row_of_pixels <= 8'b00110110;
		12'd2499: row_of_pixels <= 8'b00100110;
		12'd2500: row_of_pixels <= 8'b00000110;
		12'd2501: row_of_pixels <= 8'b00001111;
		12'd2502: row_of_pixels <= 8'b00000110;
		12'd2503: row_of_pixels <= 8'b00000110;
		12'd2504: row_of_pixels <= 8'b00000110;
		12'd2505: row_of_pixels <= 8'b00000110;
		12'd2506: row_of_pixels <= 8'b01100111;
		12'd2507: row_of_pixels <= 8'b00111111;
		12'd2508: row_of_pixels <= 8'b00000000;
		12'd2509: row_of_pixels <= 8'b00000000;
		12'd2510: row_of_pixels <= 8'b00000000;
		12'd2511: row_of_pixels <= 8'b00000000;
		12'd2512: row_of_pixels <= 8'b00000000;
		12'd2513: row_of_pixels <= 8'b00000000;
		12'd2514: row_of_pixels <= 8'b11000011;
		12'd2515: row_of_pixels <= 8'b01100110;
		12'd2516: row_of_pixels <= 8'b00111100;
		12'd2517: row_of_pixels <= 8'b00011000;
		12'd2518: row_of_pixels <= 8'b11111111;
		12'd2519: row_of_pixels <= 8'b00011000;
		12'd2520: row_of_pixels <= 8'b11111111;
		12'd2521: row_of_pixels <= 8'b00011000;
		12'd2522: row_of_pixels <= 8'b00011000;
		12'd2523: row_of_pixels <= 8'b00011000;
		12'd2524: row_of_pixels <= 8'b00000000;
		12'd2525: row_of_pixels <= 8'b00000000;
		12'd2526: row_of_pixels <= 8'b00000000;
		12'd2527: row_of_pixels <= 8'b00000000;
		12'd2528: row_of_pixels <= 8'b00000000;
		12'd2529: row_of_pixels <= 8'b00111111;
		12'd2530: row_of_pixels <= 8'b01100110;
		12'd2531: row_of_pixels <= 8'b01100110;
		12'd2532: row_of_pixels <= 8'b00111110;
		12'd2533: row_of_pixels <= 8'b01000110;
		12'd2534: row_of_pixels <= 8'b01100110;
		12'd2535: row_of_pixels <= 8'b11110110;
		12'd2536: row_of_pixels <= 8'b01100110;
		12'd2537: row_of_pixels <= 8'b01100110;
		12'd2538: row_of_pixels <= 8'b01100110;
		12'd2539: row_of_pixels <= 8'b11001111;
		12'd2540: row_of_pixels <= 8'b00000000;
		12'd2541: row_of_pixels <= 8'b00000000;
		12'd2542: row_of_pixels <= 8'b00000000;
		12'd2543: row_of_pixels <= 8'b00000000;
		12'd2544: row_of_pixels <= 8'b00000000;
		12'd2545: row_of_pixels <= 8'b01110000;
		12'd2546: row_of_pixels <= 8'b11011000;
		12'd2547: row_of_pixels <= 8'b00011000;
		12'd2548: row_of_pixels <= 8'b00011000;
		12'd2549: row_of_pixels <= 8'b00011000;
		12'd2550: row_of_pixels <= 8'b01111110;
		12'd2551: row_of_pixels <= 8'b00011000;
		12'd2552: row_of_pixels <= 8'b00011000;
		12'd2553: row_of_pixels <= 8'b00011000;
		12'd2554: row_of_pixels <= 8'b00011000;
		12'd2555: row_of_pixels <= 8'b00011000;
		12'd2556: row_of_pixels <= 8'b00011011;
		12'd2557: row_of_pixels <= 8'b00001110;
		12'd2558: row_of_pixels <= 8'b00000000;
		12'd2559: row_of_pixels <= 8'b00000000;
		12'd2560: row_of_pixels <= 8'b00000000;
		12'd2561: row_of_pixels <= 8'b00011000;
		12'd2562: row_of_pixels <= 8'b00001100;
		12'd2563: row_of_pixels <= 8'b00000110;
		12'd2564: row_of_pixels <= 8'b00000000;
		12'd2565: row_of_pixels <= 8'b00011110;
		12'd2566: row_of_pixels <= 8'b00110000;
		12'd2567: row_of_pixels <= 8'b00111110;
		12'd2568: row_of_pixels <= 8'b00110011;
		12'd2569: row_of_pixels <= 8'b00110011;
		12'd2570: row_of_pixels <= 8'b00110011;
		12'd2571: row_of_pixels <= 8'b01101110;
		12'd2572: row_of_pixels <= 8'b00000000;
		12'd2573: row_of_pixels <= 8'b00000000;
		12'd2574: row_of_pixels <= 8'b00000000;
		12'd2575: row_of_pixels <= 8'b00000000;
		12'd2576: row_of_pixels <= 8'b00000000;
		12'd2577: row_of_pixels <= 8'b00110000;
		12'd2578: row_of_pixels <= 8'b00011000;
		12'd2579: row_of_pixels <= 8'b00001100;
		12'd2580: row_of_pixels <= 8'b00000000;
		12'd2581: row_of_pixels <= 8'b00011100;
		12'd2582: row_of_pixels <= 8'b00011000;
		12'd2583: row_of_pixels <= 8'b00011000;
		12'd2584: row_of_pixels <= 8'b00011000;
		12'd2585: row_of_pixels <= 8'b00011000;
		12'd2586: row_of_pixels <= 8'b00011000;
		12'd2587: row_of_pixels <= 8'b00111100;
		12'd2588: row_of_pixels <= 8'b00000000;
		12'd2589: row_of_pixels <= 8'b00000000;
		12'd2590: row_of_pixels <= 8'b00000000;
		12'd2591: row_of_pixels <= 8'b00000000;
		12'd2592: row_of_pixels <= 8'b00000000;
		12'd2593: row_of_pixels <= 8'b00011000;
		12'd2594: row_of_pixels <= 8'b00001100;
		12'd2595: row_of_pixels <= 8'b00000110;
		12'd2596: row_of_pixels <= 8'b00000000;
		12'd2597: row_of_pixels <= 8'b00111110;
		12'd2598: row_of_pixels <= 8'b01100011;
		12'd2599: row_of_pixels <= 8'b01100011;
		12'd2600: row_of_pixels <= 8'b01100011;
		12'd2601: row_of_pixels <= 8'b01100011;
		12'd2602: row_of_pixels <= 8'b01100011;
		12'd2603: row_of_pixels <= 8'b00111110;
		12'd2604: row_of_pixels <= 8'b00000000;
		12'd2605: row_of_pixels <= 8'b00000000;
		12'd2606: row_of_pixels <= 8'b00000000;
		12'd2607: row_of_pixels <= 8'b00000000;
		12'd2608: row_of_pixels <= 8'b00000000;
		12'd2609: row_of_pixels <= 8'b00011000;
		12'd2610: row_of_pixels <= 8'b00001100;
		12'd2611: row_of_pixels <= 8'b00000110;
		12'd2612: row_of_pixels <= 8'b00000000;
		12'd2613: row_of_pixels <= 8'b00110011;
		12'd2614: row_of_pixels <= 8'b00110011;
		12'd2615: row_of_pixels <= 8'b00110011;
		12'd2616: row_of_pixels <= 8'b00110011;
		12'd2617: row_of_pixels <= 8'b00110011;
		12'd2618: row_of_pixels <= 8'b00110011;
		12'd2619: row_of_pixels <= 8'b01101110;
		12'd2620: row_of_pixels <= 8'b00000000;
		12'd2621: row_of_pixels <= 8'b00000000;
		12'd2622: row_of_pixels <= 8'b00000000;
		12'd2623: row_of_pixels <= 8'b00000000;
		12'd2624: row_of_pixels <= 8'b00000000;
		12'd2625: row_of_pixels <= 8'b00000000;
		12'd2626: row_of_pixels <= 8'b01101110;
		12'd2627: row_of_pixels <= 8'b00111011;
		12'd2628: row_of_pixels <= 8'b00000000;
		12'd2629: row_of_pixels <= 8'b00111011;
		12'd2630: row_of_pixels <= 8'b01100110;
		12'd2631: row_of_pixels <= 8'b01100110;
		12'd2632: row_of_pixels <= 8'b01100110;
		12'd2633: row_of_pixels <= 8'b01100110;
		12'd2634: row_of_pixels <= 8'b01100110;
		12'd2635: row_of_pixels <= 8'b01100110;
		12'd2636: row_of_pixels <= 8'b00000000;
		12'd2637: row_of_pixels <= 8'b00000000;
		12'd2638: row_of_pixels <= 8'b00000000;
		12'd2639: row_of_pixels <= 8'b00000000;
		12'd2640: row_of_pixels <= 8'b01101110;
		12'd2641: row_of_pixels <= 8'b00111011;
		12'd2642: row_of_pixels <= 8'b00000000;
		12'd2643: row_of_pixels <= 8'b01100011;
		12'd2644: row_of_pixels <= 8'b01100111;
		12'd2645: row_of_pixels <= 8'b01101111;
		12'd2646: row_of_pixels <= 8'b01111111;
		12'd2647: row_of_pixels <= 8'b01111011;
		12'd2648: row_of_pixels <= 8'b01110011;
		12'd2649: row_of_pixels <= 8'b01100011;
		12'd2650: row_of_pixels <= 8'b01100011;
		12'd2651: row_of_pixels <= 8'b01100011;
		12'd2652: row_of_pixels <= 8'b00000000;
		12'd2653: row_of_pixels <= 8'b00000000;
		12'd2654: row_of_pixels <= 8'b00000000;
		12'd2655: row_of_pixels <= 8'b00000000;
		12'd2656: row_of_pixels <= 8'b00000000;
		12'd2657: row_of_pixels <= 8'b00111100;
		12'd2658: row_of_pixels <= 8'b00110110;
		12'd2659: row_of_pixels <= 8'b00110110;
		12'd2660: row_of_pixels <= 8'b01111100;
		12'd2661: row_of_pixels <= 8'b00000000;
		12'd2662: row_of_pixels <= 8'b01111110;
		12'd2663: row_of_pixels <= 8'b00000000;
		12'd2664: row_of_pixels <= 8'b00000000;
		12'd2665: row_of_pixels <= 8'b00000000;
		12'd2666: row_of_pixels <= 8'b00000000;
		12'd2667: row_of_pixels <= 8'b00000000;
		12'd2668: row_of_pixels <= 8'b00000000;
		12'd2669: row_of_pixels <= 8'b00000000;
		12'd2670: row_of_pixels <= 8'b00000000;
		12'd2671: row_of_pixels <= 8'b00000000;
		12'd2672: row_of_pixels <= 8'b00000000;
		12'd2673: row_of_pixels <= 8'b00011100;
		12'd2674: row_of_pixels <= 8'b00110110;
		12'd2675: row_of_pixels <= 8'b00110110;
		12'd2676: row_of_pixels <= 8'b00011100;
		12'd2677: row_of_pixels <= 8'b00000000;
		12'd2678: row_of_pixels <= 8'b00111110;
		12'd2679: row_of_pixels <= 8'b00000000;
		12'd2680: row_of_pixels <= 8'b00000000;
		12'd2681: row_of_pixels <= 8'b00000000;
		12'd2682: row_of_pixels <= 8'b00000000;
		12'd2683: row_of_pixels <= 8'b00000000;
		12'd2684: row_of_pixels <= 8'b00000000;
		12'd2685: row_of_pixels <= 8'b00000000;
		12'd2686: row_of_pixels <= 8'b00000000;
		12'd2687: row_of_pixels <= 8'b00000000;
		12'd2688: row_of_pixels <= 8'b00000000;
		12'd2689: row_of_pixels <= 8'b00000000;
		12'd2690: row_of_pixels <= 8'b00001100;
		12'd2691: row_of_pixels <= 8'b00001100;
		12'd2692: row_of_pixels <= 8'b00000000;
		12'd2693: row_of_pixels <= 8'b00001100;
		12'd2694: row_of_pixels <= 8'b00001100;
		12'd2695: row_of_pixels <= 8'b00000110;
		12'd2696: row_of_pixels <= 8'b00000011;
		12'd2697: row_of_pixels <= 8'b01100011;
		12'd2698: row_of_pixels <= 8'b01100011;
		12'd2699: row_of_pixels <= 8'b00111110;
		12'd2700: row_of_pixels <= 8'b00000000;
		12'd2701: row_of_pixels <= 8'b00000000;
		12'd2702: row_of_pixels <= 8'b00000000;
		12'd2703: row_of_pixels <= 8'b00000000;
		12'd2704: row_of_pixels <= 8'b00000000;
		12'd2705: row_of_pixels <= 8'b00000000;
		12'd2706: row_of_pixels <= 8'b00000000;
		12'd2707: row_of_pixels <= 8'b00000000;
		12'd2708: row_of_pixels <= 8'b00000000;
		12'd2709: row_of_pixels <= 8'b00000000;
		12'd2710: row_of_pixels <= 8'b01111111;
		12'd2711: row_of_pixels <= 8'b00000011;
		12'd2712: row_of_pixels <= 8'b00000011;
		12'd2713: row_of_pixels <= 8'b00000011;
		12'd2714: row_of_pixels <= 8'b00000011;
		12'd2715: row_of_pixels <= 8'b00000000;
		12'd2716: row_of_pixels <= 8'b00000000;
		12'd2717: row_of_pixels <= 8'b00000000;
		12'd2718: row_of_pixels <= 8'b00000000;
		12'd2719: row_of_pixels <= 8'b00000000;
		12'd2720: row_of_pixels <= 8'b00000000;
		12'd2721: row_of_pixels <= 8'b00000000;
		12'd2722: row_of_pixels <= 8'b00000000;
		12'd2723: row_of_pixels <= 8'b00000000;
		12'd2724: row_of_pixels <= 8'b00000000;
		12'd2725: row_of_pixels <= 8'b00000000;
		12'd2726: row_of_pixels <= 8'b01111111;
		12'd2727: row_of_pixels <= 8'b01100000;
		12'd2728: row_of_pixels <= 8'b01100000;
		12'd2729: row_of_pixels <= 8'b01100000;
		12'd2730: row_of_pixels <= 8'b01100000;
		12'd2731: row_of_pixels <= 8'b00000000;
		12'd2732: row_of_pixels <= 8'b00000000;
		12'd2733: row_of_pixels <= 8'b00000000;
		12'd2734: row_of_pixels <= 8'b00000000;
		12'd2735: row_of_pixels <= 8'b00000000;
		12'd2736: row_of_pixels <= 8'b00000000;
		12'd2737: row_of_pixels <= 8'b00000011;
		12'd2738: row_of_pixels <= 8'b00000011;
		12'd2739: row_of_pixels <= 8'b01000011;
		12'd2740: row_of_pixels <= 8'b01100011;
		12'd2741: row_of_pixels <= 8'b00110011;
		12'd2742: row_of_pixels <= 8'b00011000;
		12'd2743: row_of_pixels <= 8'b00001100;
		12'd2744: row_of_pixels <= 8'b00000110;
		12'd2745: row_of_pixels <= 8'b01110011;
		12'd2746: row_of_pixels <= 8'b11011001;
		12'd2747: row_of_pixels <= 8'b01100000;
		12'd2748: row_of_pixels <= 8'b00110000;
		12'd2749: row_of_pixels <= 8'b11111000;
		12'd2750: row_of_pixels <= 8'b00000000;
		12'd2751: row_of_pixels <= 8'b00000000;
		12'd2752: row_of_pixels <= 8'b00000000;
		12'd2753: row_of_pixels <= 8'b00000011;
		12'd2754: row_of_pixels <= 8'b00000011;
		12'd2755: row_of_pixels <= 8'b01000011;
		12'd2756: row_of_pixels <= 8'b01100011;
		12'd2757: row_of_pixels <= 8'b00110011;
		12'd2758: row_of_pixels <= 8'b00011000;
		12'd2759: row_of_pixels <= 8'b00001100;
		12'd2760: row_of_pixels <= 8'b01100110;
		12'd2761: row_of_pixels <= 8'b01110011;
		12'd2762: row_of_pixels <= 8'b01101001;
		12'd2763: row_of_pixels <= 8'b01111100;
		12'd2764: row_of_pixels <= 8'b01100000;
		12'd2765: row_of_pixels <= 8'b01100000;
		12'd2766: row_of_pixels <= 8'b00000000;
		12'd2767: row_of_pixels <= 8'b00000000;
		12'd2768: row_of_pixels <= 8'b00000000;
		12'd2769: row_of_pixels <= 8'b00000000;
		12'd2770: row_of_pixels <= 8'b00011000;
		12'd2771: row_of_pixels <= 8'b00011000;
		12'd2772: row_of_pixels <= 8'b00000000;
		12'd2773: row_of_pixels <= 8'b00011000;
		12'd2774: row_of_pixels <= 8'b00011000;
		12'd2775: row_of_pixels <= 8'b00011000;
		12'd2776: row_of_pixels <= 8'b00111100;
		12'd2777: row_of_pixels <= 8'b00111100;
		12'd2778: row_of_pixels <= 8'b00111100;
		12'd2779: row_of_pixels <= 8'b00011000;
		12'd2780: row_of_pixels <= 8'b00000000;
		12'd2781: row_of_pixels <= 8'b00000000;
		12'd2782: row_of_pixels <= 8'b00000000;
		12'd2783: row_of_pixels <= 8'b00000000;
		12'd2784: row_of_pixels <= 8'b00000000;
		12'd2785: row_of_pixels <= 8'b00000000;
		12'd2786: row_of_pixels <= 8'b00000000;
		12'd2787: row_of_pixels <= 8'b00000000;
		12'd2788: row_of_pixels <= 8'b00000000;
		12'd2789: row_of_pixels <= 8'b01101100;
		12'd2790: row_of_pixels <= 8'b00110110;
		12'd2791: row_of_pixels <= 8'b00011011;
		12'd2792: row_of_pixels <= 8'b00110110;
		12'd2793: row_of_pixels <= 8'b01101100;
		12'd2794: row_of_pixels <= 8'b00000000;
		12'd2795: row_of_pixels <= 8'b00000000;
		12'd2796: row_of_pixels <= 8'b00000000;
		12'd2797: row_of_pixels <= 8'b00000000;
		12'd2798: row_of_pixels <= 8'b00000000;
		12'd2799: row_of_pixels <= 8'b00000000;
		12'd2800: row_of_pixels <= 8'b00000000;
		12'd2801: row_of_pixels <= 8'b00000000;
		12'd2802: row_of_pixels <= 8'b00000000;
		12'd2803: row_of_pixels <= 8'b00000000;
		12'd2804: row_of_pixels <= 8'b00000000;
		12'd2805: row_of_pixels <= 8'b00011011;
		12'd2806: row_of_pixels <= 8'b00110110;
		12'd2807: row_of_pixels <= 8'b01101100;
		12'd2808: row_of_pixels <= 8'b00110110;
		12'd2809: row_of_pixels <= 8'b00011011;
		12'd2810: row_of_pixels <= 8'b00000000;
		12'd2811: row_of_pixels <= 8'b00000000;
		12'd2812: row_of_pixels <= 8'b00000000;
		12'd2813: row_of_pixels <= 8'b00000000;
		12'd2814: row_of_pixels <= 8'b00000000;
		12'd2815: row_of_pixels <= 8'b00000000;
		12'd2816: row_of_pixels <= 8'b10001000;
		12'd2817: row_of_pixels <= 8'b00100010;
		12'd2818: row_of_pixels <= 8'b10001000;
		12'd2819: row_of_pixels <= 8'b00100010;
		12'd2820: row_of_pixels <= 8'b10001000;
		12'd2821: row_of_pixels <= 8'b00100010;
		12'd2822: row_of_pixels <= 8'b10001000;
		12'd2823: row_of_pixels <= 8'b00100010;
		12'd2824: row_of_pixels <= 8'b10001000;
		12'd2825: row_of_pixels <= 8'b00100010;
		12'd2826: row_of_pixels <= 8'b10001000;
		12'd2827: row_of_pixels <= 8'b00100010;
		12'd2828: row_of_pixels <= 8'b10001000;
		12'd2829: row_of_pixels <= 8'b00100010;
		12'd2830: row_of_pixels <= 8'b10001000;
		12'd2831: row_of_pixels <= 8'b00100010;
		12'd2832: row_of_pixels <= 8'b10101010;
		12'd2833: row_of_pixels <= 8'b01010101;
		12'd2834: row_of_pixels <= 8'b10101010;
		12'd2835: row_of_pixels <= 8'b01010101;
		12'd2836: row_of_pixels <= 8'b10101010;
		12'd2837: row_of_pixels <= 8'b01010101;
		12'd2838: row_of_pixels <= 8'b10101010;
		12'd2839: row_of_pixels <= 8'b01010101;
		12'd2840: row_of_pixels <= 8'b10101010;
		12'd2841: row_of_pixels <= 8'b01010101;
		12'd2842: row_of_pixels <= 8'b10101010;
		12'd2843: row_of_pixels <= 8'b01010101;
		12'd2844: row_of_pixels <= 8'b10101010;
		12'd2845: row_of_pixels <= 8'b01010101;
		12'd2846: row_of_pixels <= 8'b10101010;
		12'd2847: row_of_pixels <= 8'b01010101;
		12'd2848: row_of_pixels <= 8'b10111011;
		12'd2849: row_of_pixels <= 8'b11101110;
		12'd2850: row_of_pixels <= 8'b10111011;
		12'd2851: row_of_pixels <= 8'b11101110;
		12'd2852: row_of_pixels <= 8'b10111011;
		12'd2853: row_of_pixels <= 8'b11101110;
		12'd2854: row_of_pixels <= 8'b10111011;
		12'd2855: row_of_pixels <= 8'b11101110;
		12'd2856: row_of_pixels <= 8'b10111011;
		12'd2857: row_of_pixels <= 8'b11101110;
		12'd2858: row_of_pixels <= 8'b10111011;
		12'd2859: row_of_pixels <= 8'b11101110;
		12'd2860: row_of_pixels <= 8'b10111011;
		12'd2861: row_of_pixels <= 8'b11101110;
		12'd2862: row_of_pixels <= 8'b10111011;
		12'd2863: row_of_pixels <= 8'b11101110;
		12'd2864: row_of_pixels <= 8'b00011000;
		12'd2865: row_of_pixels <= 8'b00011000;
		12'd2866: row_of_pixels <= 8'b00011000;
		12'd2867: row_of_pixels <= 8'b00011000;
		12'd2868: row_of_pixels <= 8'b00011000;
		12'd2869: row_of_pixels <= 8'b00011000;
		12'd2870: row_of_pixels <= 8'b00011000;
		12'd2871: row_of_pixels <= 8'b00011000;
		12'd2872: row_of_pixels <= 8'b00011000;
		12'd2873: row_of_pixels <= 8'b00011000;
		12'd2874: row_of_pixels <= 8'b00011000;
		12'd2875: row_of_pixels <= 8'b00011000;
		12'd2876: row_of_pixels <= 8'b00011000;
		12'd2877: row_of_pixels <= 8'b00011000;
		12'd2878: row_of_pixels <= 8'b00011000;
		12'd2879: row_of_pixels <= 8'b00011000;
		12'd2880: row_of_pixels <= 8'b00011000;
		12'd2881: row_of_pixels <= 8'b00011000;
		12'd2882: row_of_pixels <= 8'b00011000;
		12'd2883: row_of_pixels <= 8'b00011000;
		12'd2884: row_of_pixels <= 8'b00011000;
		12'd2885: row_of_pixels <= 8'b00011000;
		12'd2886: row_of_pixels <= 8'b00011000;
		12'd2887: row_of_pixels <= 8'b00011111;
		12'd2888: row_of_pixels <= 8'b00011000;
		12'd2889: row_of_pixels <= 8'b00011000;
		12'd2890: row_of_pixels <= 8'b00011000;
		12'd2891: row_of_pixels <= 8'b00011000;
		12'd2892: row_of_pixels <= 8'b00011000;
		12'd2893: row_of_pixels <= 8'b00011000;
		12'd2894: row_of_pixels <= 8'b00011000;
		12'd2895: row_of_pixels <= 8'b00011000;
		12'd2896: row_of_pixels <= 8'b00011000;
		12'd2897: row_of_pixels <= 8'b00011000;
		12'd2898: row_of_pixels <= 8'b00011000;
		12'd2899: row_of_pixels <= 8'b00011000;
		12'd2900: row_of_pixels <= 8'b00011000;
		12'd2901: row_of_pixels <= 8'b00011111;
		12'd2902: row_of_pixels <= 8'b00011000;
		12'd2903: row_of_pixels <= 8'b00011111;
		12'd2904: row_of_pixels <= 8'b00011000;
		12'd2905: row_of_pixels <= 8'b00011000;
		12'd2906: row_of_pixels <= 8'b00011000;
		12'd2907: row_of_pixels <= 8'b00011000;
		12'd2908: row_of_pixels <= 8'b00011000;
		12'd2909: row_of_pixels <= 8'b00011000;
		12'd2910: row_of_pixels <= 8'b00011000;
		12'd2911: row_of_pixels <= 8'b00011000;
		12'd2912: row_of_pixels <= 8'b01101100;
		12'd2913: row_of_pixels <= 8'b01101100;
		12'd2914: row_of_pixels <= 8'b01101100;
		12'd2915: row_of_pixels <= 8'b01101100;
		12'd2916: row_of_pixels <= 8'b01101100;
		12'd2917: row_of_pixels <= 8'b01101100;
		12'd2918: row_of_pixels <= 8'b01101100;
		12'd2919: row_of_pixels <= 8'b01101111;
		12'd2920: row_of_pixels <= 8'b01101100;
		12'd2921: row_of_pixels <= 8'b01101100;
		12'd2922: row_of_pixels <= 8'b01101100;
		12'd2923: row_of_pixels <= 8'b01101100;
		12'd2924: row_of_pixels <= 8'b01101100;
		12'd2925: row_of_pixels <= 8'b01101100;
		12'd2926: row_of_pixels <= 8'b01101100;
		12'd2927: row_of_pixels <= 8'b01101100;
		12'd2928: row_of_pixels <= 8'b00000000;
		12'd2929: row_of_pixels <= 8'b00000000;
		12'd2930: row_of_pixels <= 8'b00000000;
		12'd2931: row_of_pixels <= 8'b00000000;
		12'd2932: row_of_pixels <= 8'b00000000;
		12'd2933: row_of_pixels <= 8'b00000000;
		12'd2934: row_of_pixels <= 8'b00000000;
		12'd2935: row_of_pixels <= 8'b01111111;
		12'd2936: row_of_pixels <= 8'b01101100;
		12'd2937: row_of_pixels <= 8'b01101100;
		12'd2938: row_of_pixels <= 8'b01101100;
		12'd2939: row_of_pixels <= 8'b01101100;
		12'd2940: row_of_pixels <= 8'b01101100;
		12'd2941: row_of_pixels <= 8'b01101100;
		12'd2942: row_of_pixels <= 8'b01101100;
		12'd2943: row_of_pixels <= 8'b01101100;
		12'd2944: row_of_pixels <= 8'b00000000;
		12'd2945: row_of_pixels <= 8'b00000000;
		12'd2946: row_of_pixels <= 8'b00000000;
		12'd2947: row_of_pixels <= 8'b00000000;
		12'd2948: row_of_pixels <= 8'b00000000;
		12'd2949: row_of_pixels <= 8'b00011111;
		12'd2950: row_of_pixels <= 8'b00011000;
		12'd2951: row_of_pixels <= 8'b00011111;
		12'd2952: row_of_pixels <= 8'b00011000;
		12'd2953: row_of_pixels <= 8'b00011000;
		12'd2954: row_of_pixels <= 8'b00011000;
		12'd2955: row_of_pixels <= 8'b00011000;
		12'd2956: row_of_pixels <= 8'b00011000;
		12'd2957: row_of_pixels <= 8'b00011000;
		12'd2958: row_of_pixels <= 8'b00011000;
		12'd2959: row_of_pixels <= 8'b00011000;
		12'd2960: row_of_pixels <= 8'b01101100;
		12'd2961: row_of_pixels <= 8'b01101100;
		12'd2962: row_of_pixels <= 8'b01101100;
		12'd2963: row_of_pixels <= 8'b01101100;
		12'd2964: row_of_pixels <= 8'b01101100;
		12'd2965: row_of_pixels <= 8'b01101111;
		12'd2966: row_of_pixels <= 8'b01100000;
		12'd2967: row_of_pixels <= 8'b01101111;
		12'd2968: row_of_pixels <= 8'b01101100;
		12'd2969: row_of_pixels <= 8'b01101100;
		12'd2970: row_of_pixels <= 8'b01101100;
		12'd2971: row_of_pixels <= 8'b01101100;
		12'd2972: row_of_pixels <= 8'b01101100;
		12'd2973: row_of_pixels <= 8'b01101100;
		12'd2974: row_of_pixels <= 8'b01101100;
		12'd2975: row_of_pixels <= 8'b01101100;
		12'd2976: row_of_pixels <= 8'b01101100;
		12'd2977: row_of_pixels <= 8'b01101100;
		12'd2978: row_of_pixels <= 8'b01101100;
		12'd2979: row_of_pixels <= 8'b01101100;
		12'd2980: row_of_pixels <= 8'b01101100;
		12'd2981: row_of_pixels <= 8'b01101100;
		12'd2982: row_of_pixels <= 8'b01101100;
		12'd2983: row_of_pixels <= 8'b01101100;
		12'd2984: row_of_pixels <= 8'b01101100;
		12'd2985: row_of_pixels <= 8'b01101100;
		12'd2986: row_of_pixels <= 8'b01101100;
		12'd2987: row_of_pixels <= 8'b01101100;
		12'd2988: row_of_pixels <= 8'b01101100;
		12'd2989: row_of_pixels <= 8'b01101100;
		12'd2990: row_of_pixels <= 8'b01101100;
		12'd2991: row_of_pixels <= 8'b01101100;
		12'd2992: row_of_pixels <= 8'b00000000;
		12'd2993: row_of_pixels <= 8'b00000000;
		12'd2994: row_of_pixels <= 8'b00000000;
		12'd2995: row_of_pixels <= 8'b00000000;
		12'd2996: row_of_pixels <= 8'b00000000;
		12'd2997: row_of_pixels <= 8'b01111111;
		12'd2998: row_of_pixels <= 8'b01100000;
		12'd2999: row_of_pixels <= 8'b01101111;
		12'd3000: row_of_pixels <= 8'b01101100;
		12'd3001: row_of_pixels <= 8'b01101100;
		12'd3002: row_of_pixels <= 8'b01101100;
		12'd3003: row_of_pixels <= 8'b01101100;
		12'd3004: row_of_pixels <= 8'b01101100;
		12'd3005: row_of_pixels <= 8'b01101100;
		12'd3006: row_of_pixels <= 8'b01101100;
		12'd3007: row_of_pixels <= 8'b01101100;
		12'd3008: row_of_pixels <= 8'b01101100;
		12'd3009: row_of_pixels <= 8'b01101100;
		12'd3010: row_of_pixels <= 8'b01101100;
		12'd3011: row_of_pixels <= 8'b01101100;
		12'd3012: row_of_pixels <= 8'b01101100;
		12'd3013: row_of_pixels <= 8'b01101111;
		12'd3014: row_of_pixels <= 8'b01100000;
		12'd3015: row_of_pixels <= 8'b01111111;
		12'd3016: row_of_pixels <= 8'b00000000;
		12'd3017: row_of_pixels <= 8'b00000000;
		12'd3018: row_of_pixels <= 8'b00000000;
		12'd3019: row_of_pixels <= 8'b00000000;
		12'd3020: row_of_pixels <= 8'b00000000;
		12'd3021: row_of_pixels <= 8'b00000000;
		12'd3022: row_of_pixels <= 8'b00000000;
		12'd3023: row_of_pixels <= 8'b00000000;
		12'd3024: row_of_pixels <= 8'b01101100;
		12'd3025: row_of_pixels <= 8'b01101100;
		12'd3026: row_of_pixels <= 8'b01101100;
		12'd3027: row_of_pixels <= 8'b01101100;
		12'd3028: row_of_pixels <= 8'b01101100;
		12'd3029: row_of_pixels <= 8'b01101100;
		12'd3030: row_of_pixels <= 8'b01101100;
		12'd3031: row_of_pixels <= 8'b01111111;
		12'd3032: row_of_pixels <= 8'b00000000;
		12'd3033: row_of_pixels <= 8'b00000000;
		12'd3034: row_of_pixels <= 8'b00000000;
		12'd3035: row_of_pixels <= 8'b00000000;
		12'd3036: row_of_pixels <= 8'b00000000;
		12'd3037: row_of_pixels <= 8'b00000000;
		12'd3038: row_of_pixels <= 8'b00000000;
		12'd3039: row_of_pixels <= 8'b00000000;
		12'd3040: row_of_pixels <= 8'b00011000;
		12'd3041: row_of_pixels <= 8'b00011000;
		12'd3042: row_of_pixels <= 8'b00011000;
		12'd3043: row_of_pixels <= 8'b00011000;
		12'd3044: row_of_pixels <= 8'b00011000;
		12'd3045: row_of_pixels <= 8'b00011111;
		12'd3046: row_of_pixels <= 8'b00011000;
		12'd3047: row_of_pixels <= 8'b00011111;
		12'd3048: row_of_pixels <= 8'b00000000;
		12'd3049: row_of_pixels <= 8'b00000000;
		12'd3050: row_of_pixels <= 8'b00000000;
		12'd3051: row_of_pixels <= 8'b00000000;
		12'd3052: row_of_pixels <= 8'b00000000;
		12'd3053: row_of_pixels <= 8'b00000000;
		12'd3054: row_of_pixels <= 8'b00000000;
		12'd3055: row_of_pixels <= 8'b00000000;
		12'd3056: row_of_pixels <= 8'b00000000;
		12'd3057: row_of_pixels <= 8'b00000000;
		12'd3058: row_of_pixels <= 8'b00000000;
		12'd3059: row_of_pixels <= 8'b00000000;
		12'd3060: row_of_pixels <= 8'b00000000;
		12'd3061: row_of_pixels <= 8'b00000000;
		12'd3062: row_of_pixels <= 8'b00000000;
		12'd3063: row_of_pixels <= 8'b00011111;
		12'd3064: row_of_pixels <= 8'b00011000;
		12'd3065: row_of_pixels <= 8'b00011000;
		12'd3066: row_of_pixels <= 8'b00011000;
		12'd3067: row_of_pixels <= 8'b00011000;
		12'd3068: row_of_pixels <= 8'b00011000;
		12'd3069: row_of_pixels <= 8'b00011000;
		12'd3070: row_of_pixels <= 8'b00011000;
		12'd3071: row_of_pixels <= 8'b00011000;
		12'd3072: row_of_pixels <= 8'b00011000;
		12'd3073: row_of_pixels <= 8'b00011000;
		12'd3074: row_of_pixels <= 8'b00011000;
		12'd3075: row_of_pixels <= 8'b00011000;
		12'd3076: row_of_pixels <= 8'b00011000;
		12'd3077: row_of_pixels <= 8'b00011000;
		12'd3078: row_of_pixels <= 8'b00011000;
		12'd3079: row_of_pixels <= 8'b11111000;
		12'd3080: row_of_pixels <= 8'b00000000;
		12'd3081: row_of_pixels <= 8'b00000000;
		12'd3082: row_of_pixels <= 8'b00000000;
		12'd3083: row_of_pixels <= 8'b00000000;
		12'd3084: row_of_pixels <= 8'b00000000;
		12'd3085: row_of_pixels <= 8'b00000000;
		12'd3086: row_of_pixels <= 8'b00000000;
		12'd3087: row_of_pixels <= 8'b00000000;
		12'd3088: row_of_pixels <= 8'b00011000;
		12'd3089: row_of_pixels <= 8'b00011000;
		12'd3090: row_of_pixels <= 8'b00011000;
		12'd3091: row_of_pixels <= 8'b00011000;
		12'd3092: row_of_pixels <= 8'b00011000;
		12'd3093: row_of_pixels <= 8'b00011000;
		12'd3094: row_of_pixels <= 8'b00011000;
		12'd3095: row_of_pixels <= 8'b11111111;
		12'd3096: row_of_pixels <= 8'b00000000;
		12'd3097: row_of_pixels <= 8'b00000000;
		12'd3098: row_of_pixels <= 8'b00000000;
		12'd3099: row_of_pixels <= 8'b00000000;
		12'd3100: row_of_pixels <= 8'b00000000;
		12'd3101: row_of_pixels <= 8'b00000000;
		12'd3102: row_of_pixels <= 8'b00000000;
		12'd3103: row_of_pixels <= 8'b00000000;
		12'd3104: row_of_pixels <= 8'b00000000;
		12'd3105: row_of_pixels <= 8'b00000000;
		12'd3106: row_of_pixels <= 8'b00000000;
		12'd3107: row_of_pixels <= 8'b00000000;
		12'd3108: row_of_pixels <= 8'b00000000;
		12'd3109: row_of_pixels <= 8'b00000000;
		12'd3110: row_of_pixels <= 8'b00000000;
		12'd3111: row_of_pixels <= 8'b11111111;
		12'd3112: row_of_pixels <= 8'b00011000;
		12'd3113: row_of_pixels <= 8'b00011000;
		12'd3114: row_of_pixels <= 8'b00011000;
		12'd3115: row_of_pixels <= 8'b00011000;
		12'd3116: row_of_pixels <= 8'b00011000;
		12'd3117: row_of_pixels <= 8'b00011000;
		12'd3118: row_of_pixels <= 8'b00011000;
		12'd3119: row_of_pixels <= 8'b00011000;
		12'd3120: row_of_pixels <= 8'b00011000;
		12'd3121: row_of_pixels <= 8'b00011000;
		12'd3122: row_of_pixels <= 8'b00011000;
		12'd3123: row_of_pixels <= 8'b00011000;
		12'd3124: row_of_pixels <= 8'b00011000;
		12'd3125: row_of_pixels <= 8'b00011000;
		12'd3126: row_of_pixels <= 8'b00011000;
		12'd3127: row_of_pixels <= 8'b11111000;
		12'd3128: row_of_pixels <= 8'b00011000;
		12'd3129: row_of_pixels <= 8'b00011000;
		12'd3130: row_of_pixels <= 8'b00011000;
		12'd3131: row_of_pixels <= 8'b00011000;
		12'd3132: row_of_pixels <= 8'b00011000;
		12'd3133: row_of_pixels <= 8'b00011000;
		12'd3134: row_of_pixels <= 8'b00011000;
		12'd3135: row_of_pixels <= 8'b00011000;
		12'd3136: row_of_pixels <= 8'b00000000;
		12'd3137: row_of_pixels <= 8'b00000000;
		12'd3138: row_of_pixels <= 8'b00000000;
		12'd3139: row_of_pixels <= 8'b00000000;
		12'd3140: row_of_pixels <= 8'b00000000;
		12'd3141: row_of_pixels <= 8'b00000000;
		12'd3142: row_of_pixels <= 8'b00000000;
		12'd3143: row_of_pixels <= 8'b11111111;
		12'd3144: row_of_pixels <= 8'b00000000;
		12'd3145: row_of_pixels <= 8'b00000000;
		12'd3146: row_of_pixels <= 8'b00000000;
		12'd3147: row_of_pixels <= 8'b00000000;
		12'd3148: row_of_pixels <= 8'b00000000;
		12'd3149: row_of_pixels <= 8'b00000000;
		12'd3150: row_of_pixels <= 8'b00000000;
		12'd3151: row_of_pixels <= 8'b00000000;
		12'd3152: row_of_pixels <= 8'b00011000;
		12'd3153: row_of_pixels <= 8'b00011000;
		12'd3154: row_of_pixels <= 8'b00011000;
		12'd3155: row_of_pixels <= 8'b00011000;
		12'd3156: row_of_pixels <= 8'b00011000;
		12'd3157: row_of_pixels <= 8'b00011000;
		12'd3158: row_of_pixels <= 8'b00011000;
		12'd3159: row_of_pixels <= 8'b11111111;
		12'd3160: row_of_pixels <= 8'b00011000;
		12'd3161: row_of_pixels <= 8'b00011000;
		12'd3162: row_of_pixels <= 8'b00011000;
		12'd3163: row_of_pixels <= 8'b00011000;
		12'd3164: row_of_pixels <= 8'b00011000;
		12'd3165: row_of_pixels <= 8'b00011000;
		12'd3166: row_of_pixels <= 8'b00011000;
		12'd3167: row_of_pixels <= 8'b00011000;
		12'd3168: row_of_pixels <= 8'b00011000;
		12'd3169: row_of_pixels <= 8'b00011000;
		12'd3170: row_of_pixels <= 8'b00011000;
		12'd3171: row_of_pixels <= 8'b00011000;
		12'd3172: row_of_pixels <= 8'b00011000;
		12'd3173: row_of_pixels <= 8'b11111000;
		12'd3174: row_of_pixels <= 8'b00011000;
		12'd3175: row_of_pixels <= 8'b11111000;
		12'd3176: row_of_pixels <= 8'b00011000;
		12'd3177: row_of_pixels <= 8'b00011000;
		12'd3178: row_of_pixels <= 8'b00011000;
		12'd3179: row_of_pixels <= 8'b00011000;
		12'd3180: row_of_pixels <= 8'b00011000;
		12'd3181: row_of_pixels <= 8'b00011000;
		12'd3182: row_of_pixels <= 8'b00011000;
		12'd3183: row_of_pixels <= 8'b00011000;
		12'd3184: row_of_pixels <= 8'b01101100;
		12'd3185: row_of_pixels <= 8'b01101100;
		12'd3186: row_of_pixels <= 8'b01101100;
		12'd3187: row_of_pixels <= 8'b01101100;
		12'd3188: row_of_pixels <= 8'b01101100;
		12'd3189: row_of_pixels <= 8'b01101100;
		12'd3190: row_of_pixels <= 8'b01101100;
		12'd3191: row_of_pixels <= 8'b11101100;
		12'd3192: row_of_pixels <= 8'b01101100;
		12'd3193: row_of_pixels <= 8'b01101100;
		12'd3194: row_of_pixels <= 8'b01101100;
		12'd3195: row_of_pixels <= 8'b01101100;
		12'd3196: row_of_pixels <= 8'b01101100;
		12'd3197: row_of_pixels <= 8'b01101100;
		12'd3198: row_of_pixels <= 8'b01101100;
		12'd3199: row_of_pixels <= 8'b01101100;
		12'd3200: row_of_pixels <= 8'b01101100;
		12'd3201: row_of_pixels <= 8'b01101100;
		12'd3202: row_of_pixels <= 8'b01101100;
		12'd3203: row_of_pixels <= 8'b01101100;
		12'd3204: row_of_pixels <= 8'b01101100;
		12'd3205: row_of_pixels <= 8'b11101100;
		12'd3206: row_of_pixels <= 8'b00001100;
		12'd3207: row_of_pixels <= 8'b11111100;
		12'd3208: row_of_pixels <= 8'b00000000;
		12'd3209: row_of_pixels <= 8'b00000000;
		12'd3210: row_of_pixels <= 8'b00000000;
		12'd3211: row_of_pixels <= 8'b00000000;
		12'd3212: row_of_pixels <= 8'b00000000;
		12'd3213: row_of_pixels <= 8'b00000000;
		12'd3214: row_of_pixels <= 8'b00000000;
		12'd3215: row_of_pixels <= 8'b00000000;
		12'd3216: row_of_pixels <= 8'b00000000;
		12'd3217: row_of_pixels <= 8'b00000000;
		12'd3218: row_of_pixels <= 8'b00000000;
		12'd3219: row_of_pixels <= 8'b00000000;
		12'd3220: row_of_pixels <= 8'b00000000;
		12'd3221: row_of_pixels <= 8'b11111100;
		12'd3222: row_of_pixels <= 8'b00001100;
		12'd3223: row_of_pixels <= 8'b11101100;
		12'd3224: row_of_pixels <= 8'b01101100;
		12'd3225: row_of_pixels <= 8'b01101100;
		12'd3226: row_of_pixels <= 8'b01101100;
		12'd3227: row_of_pixels <= 8'b01101100;
		12'd3228: row_of_pixels <= 8'b01101100;
		12'd3229: row_of_pixels <= 8'b01101100;
		12'd3230: row_of_pixels <= 8'b01101100;
		12'd3231: row_of_pixels <= 8'b01101100;
		12'd3232: row_of_pixels <= 8'b01101100;
		12'd3233: row_of_pixels <= 8'b01101100;
		12'd3234: row_of_pixels <= 8'b01101100;
		12'd3235: row_of_pixels <= 8'b01101100;
		12'd3236: row_of_pixels <= 8'b01101100;
		12'd3237: row_of_pixels <= 8'b11101111;
		12'd3238: row_of_pixels <= 8'b00000000;
		12'd3239: row_of_pixels <= 8'b11111111;
		12'd3240: row_of_pixels <= 8'b00000000;
		12'd3241: row_of_pixels <= 8'b00000000;
		12'd3242: row_of_pixels <= 8'b00000000;
		12'd3243: row_of_pixels <= 8'b00000000;
		12'd3244: row_of_pixels <= 8'b00000000;
		12'd3245: row_of_pixels <= 8'b00000000;
		12'd3246: row_of_pixels <= 8'b00000000;
		12'd3247: row_of_pixels <= 8'b00000000;
		12'd3248: row_of_pixels <= 8'b00000000;
		12'd3249: row_of_pixels <= 8'b00000000;
		12'd3250: row_of_pixels <= 8'b00000000;
		12'd3251: row_of_pixels <= 8'b00000000;
		12'd3252: row_of_pixels <= 8'b00000000;
		12'd3253: row_of_pixels <= 8'b11111111;
		12'd3254: row_of_pixels <= 8'b00000000;
		12'd3255: row_of_pixels <= 8'b11101111;
		12'd3256: row_of_pixels <= 8'b01101100;
		12'd3257: row_of_pixels <= 8'b01101100;
		12'd3258: row_of_pixels <= 8'b01101100;
		12'd3259: row_of_pixels <= 8'b01101100;
		12'd3260: row_of_pixels <= 8'b01101100;
		12'd3261: row_of_pixels <= 8'b01101100;
		12'd3262: row_of_pixels <= 8'b01101100;
		12'd3263: row_of_pixels <= 8'b01101100;
		12'd3264: row_of_pixels <= 8'b01101100;
		12'd3265: row_of_pixels <= 8'b01101100;
		12'd3266: row_of_pixels <= 8'b01101100;
		12'd3267: row_of_pixels <= 8'b01101100;
		12'd3268: row_of_pixels <= 8'b01101100;
		12'd3269: row_of_pixels <= 8'b11101100;
		12'd3270: row_of_pixels <= 8'b00001100;
		12'd3271: row_of_pixels <= 8'b11101100;
		12'd3272: row_of_pixels <= 8'b01101100;
		12'd3273: row_of_pixels <= 8'b01101100;
		12'd3274: row_of_pixels <= 8'b01101100;
		12'd3275: row_of_pixels <= 8'b01101100;
		12'd3276: row_of_pixels <= 8'b01101100;
		12'd3277: row_of_pixels <= 8'b01101100;
		12'd3278: row_of_pixels <= 8'b01101100;
		12'd3279: row_of_pixels <= 8'b01101100;
		12'd3280: row_of_pixels <= 8'b00000000;
		12'd3281: row_of_pixels <= 8'b00000000;
		12'd3282: row_of_pixels <= 8'b00000000;
		12'd3283: row_of_pixels <= 8'b00000000;
		12'd3284: row_of_pixels <= 8'b00000000;
		12'd3285: row_of_pixels <= 8'b11111111;
		12'd3286: row_of_pixels <= 8'b00000000;
		12'd3287: row_of_pixels <= 8'b11111111;
		12'd3288: row_of_pixels <= 8'b00000000;
		12'd3289: row_of_pixels <= 8'b00000000;
		12'd3290: row_of_pixels <= 8'b00000000;
		12'd3291: row_of_pixels <= 8'b00000000;
		12'd3292: row_of_pixels <= 8'b00000000;
		12'd3293: row_of_pixels <= 8'b00000000;
		12'd3294: row_of_pixels <= 8'b00000000;
		12'd3295: row_of_pixels <= 8'b00000000;
		12'd3296: row_of_pixels <= 8'b01101100;
		12'd3297: row_of_pixels <= 8'b01101100;
		12'd3298: row_of_pixels <= 8'b01101100;
		12'd3299: row_of_pixels <= 8'b01101100;
		12'd3300: row_of_pixels <= 8'b01101100;
		12'd3301: row_of_pixels <= 8'b11101111;
		12'd3302: row_of_pixels <= 8'b00000000;
		12'd3303: row_of_pixels <= 8'b11101111;
		12'd3304: row_of_pixels <= 8'b01101100;
		12'd3305: row_of_pixels <= 8'b01101100;
		12'd3306: row_of_pixels <= 8'b01101100;
		12'd3307: row_of_pixels <= 8'b01101100;
		12'd3308: row_of_pixels <= 8'b01101100;
		12'd3309: row_of_pixels <= 8'b01101100;
		12'd3310: row_of_pixels <= 8'b01101100;
		12'd3311: row_of_pixels <= 8'b01101100;
		12'd3312: row_of_pixels <= 8'b00011000;
		12'd3313: row_of_pixels <= 8'b00011000;
		12'd3314: row_of_pixels <= 8'b00011000;
		12'd3315: row_of_pixels <= 8'b00011000;
		12'd3316: row_of_pixels <= 8'b00011000;
		12'd3317: row_of_pixels <= 8'b11111111;
		12'd3318: row_of_pixels <= 8'b00000000;
		12'd3319: row_of_pixels <= 8'b11111111;
		12'd3320: row_of_pixels <= 8'b00000000;
		12'd3321: row_of_pixels <= 8'b00000000;
		12'd3322: row_of_pixels <= 8'b00000000;
		12'd3323: row_of_pixels <= 8'b00000000;
		12'd3324: row_of_pixels <= 8'b00000000;
		12'd3325: row_of_pixels <= 8'b00000000;
		12'd3326: row_of_pixels <= 8'b00000000;
		12'd3327: row_of_pixels <= 8'b00000000;
		12'd3328: row_of_pixels <= 8'b01101100;
		12'd3329: row_of_pixels <= 8'b01101100;
		12'd3330: row_of_pixels <= 8'b01101100;
		12'd3331: row_of_pixels <= 8'b01101100;
		12'd3332: row_of_pixels <= 8'b01101100;
		12'd3333: row_of_pixels <= 8'b01101100;
		12'd3334: row_of_pixels <= 8'b01101100;
		12'd3335: row_of_pixels <= 8'b11111111;
		12'd3336: row_of_pixels <= 8'b00000000;
		12'd3337: row_of_pixels <= 8'b00000000;
		12'd3338: row_of_pixels <= 8'b00000000;
		12'd3339: row_of_pixels <= 8'b00000000;
		12'd3340: row_of_pixels <= 8'b00000000;
		12'd3341: row_of_pixels <= 8'b00000000;
		12'd3342: row_of_pixels <= 8'b00000000;
		12'd3343: row_of_pixels <= 8'b00000000;
		12'd3344: row_of_pixels <= 8'b00000000;
		12'd3345: row_of_pixels <= 8'b00000000;
		12'd3346: row_of_pixels <= 8'b00000000;
		12'd3347: row_of_pixels <= 8'b00000000;
		12'd3348: row_of_pixels <= 8'b00000000;
		12'd3349: row_of_pixels <= 8'b11111111;
		12'd3350: row_of_pixels <= 8'b00000000;
		12'd3351: row_of_pixels <= 8'b11111111;
		12'd3352: row_of_pixels <= 8'b00011000;
		12'd3353: row_of_pixels <= 8'b00011000;
		12'd3354: row_of_pixels <= 8'b00011000;
		12'd3355: row_of_pixels <= 8'b00011000;
		12'd3356: row_of_pixels <= 8'b00011000;
		12'd3357: row_of_pixels <= 8'b00011000;
		12'd3358: row_of_pixels <= 8'b00011000;
		12'd3359: row_of_pixels <= 8'b00011000;
		12'd3360: row_of_pixels <= 8'b00000000;
		12'd3361: row_of_pixels <= 8'b00000000;
		12'd3362: row_of_pixels <= 8'b00000000;
		12'd3363: row_of_pixels <= 8'b00000000;
		12'd3364: row_of_pixels <= 8'b00000000;
		12'd3365: row_of_pixels <= 8'b00000000;
		12'd3366: row_of_pixels <= 8'b00000000;
		12'd3367: row_of_pixels <= 8'b11111111;
		12'd3368: row_of_pixels <= 8'b01101100;
		12'd3369: row_of_pixels <= 8'b01101100;
		12'd3370: row_of_pixels <= 8'b01101100;
		12'd3371: row_of_pixels <= 8'b01101100;
		12'd3372: row_of_pixels <= 8'b01101100;
		12'd3373: row_of_pixels <= 8'b01101100;
		12'd3374: row_of_pixels <= 8'b01101100;
		12'd3375: row_of_pixels <= 8'b01101100;
		12'd3376: row_of_pixels <= 8'b01101100;
		12'd3377: row_of_pixels <= 8'b01101100;
		12'd3378: row_of_pixels <= 8'b01101100;
		12'd3379: row_of_pixels <= 8'b01101100;
		12'd3380: row_of_pixels <= 8'b01101100;
		12'd3381: row_of_pixels <= 8'b01101100;
		12'd3382: row_of_pixels <= 8'b01101100;
		12'd3383: row_of_pixels <= 8'b11111100;
		12'd3384: row_of_pixels <= 8'b00000000;
		12'd3385: row_of_pixels <= 8'b00000000;
		12'd3386: row_of_pixels <= 8'b00000000;
		12'd3387: row_of_pixels <= 8'b00000000;
		12'd3388: row_of_pixels <= 8'b00000000;
		12'd3389: row_of_pixels <= 8'b00000000;
		12'd3390: row_of_pixels <= 8'b00000000;
		12'd3391: row_of_pixels <= 8'b00000000;
		12'd3392: row_of_pixels <= 8'b00011000;
		12'd3393: row_of_pixels <= 8'b00011000;
		12'd3394: row_of_pixels <= 8'b00011000;
		12'd3395: row_of_pixels <= 8'b00011000;
		12'd3396: row_of_pixels <= 8'b00011000;
		12'd3397: row_of_pixels <= 8'b11111000;
		12'd3398: row_of_pixels <= 8'b00011000;
		12'd3399: row_of_pixels <= 8'b11111000;
		12'd3400: row_of_pixels <= 8'b00000000;
		12'd3401: row_of_pixels <= 8'b00000000;
		12'd3402: row_of_pixels <= 8'b00000000;
		12'd3403: row_of_pixels <= 8'b00000000;
		12'd3404: row_of_pixels <= 8'b00000000;
		12'd3405: row_of_pixels <= 8'b00000000;
		12'd3406: row_of_pixels <= 8'b00000000;
		12'd3407: row_of_pixels <= 8'b00000000;
		12'd3408: row_of_pixels <= 8'b00000000;
		12'd3409: row_of_pixels <= 8'b00000000;
		12'd3410: row_of_pixels <= 8'b00000000;
		12'd3411: row_of_pixels <= 8'b00000000;
		12'd3412: row_of_pixels <= 8'b00000000;
		12'd3413: row_of_pixels <= 8'b11111000;
		12'd3414: row_of_pixels <= 8'b00011000;
		12'd3415: row_of_pixels <= 8'b11111000;
		12'd3416: row_of_pixels <= 8'b00011000;
		12'd3417: row_of_pixels <= 8'b00011000;
		12'd3418: row_of_pixels <= 8'b00011000;
		12'd3419: row_of_pixels <= 8'b00011000;
		12'd3420: row_of_pixels <= 8'b00011000;
		12'd3421: row_of_pixels <= 8'b00011000;
		12'd3422: row_of_pixels <= 8'b00011000;
		12'd3423: row_of_pixels <= 8'b00011000;
		12'd3424: row_of_pixels <= 8'b00000000;
		12'd3425: row_of_pixels <= 8'b00000000;
		12'd3426: row_of_pixels <= 8'b00000000;
		12'd3427: row_of_pixels <= 8'b00000000;
		12'd3428: row_of_pixels <= 8'b00000000;
		12'd3429: row_of_pixels <= 8'b00000000;
		12'd3430: row_of_pixels <= 8'b00000000;
		12'd3431: row_of_pixels <= 8'b11111100;
		12'd3432: row_of_pixels <= 8'b01101100;
		12'd3433: row_of_pixels <= 8'b01101100;
		12'd3434: row_of_pixels <= 8'b01101100;
		12'd3435: row_of_pixels <= 8'b01101100;
		12'd3436: row_of_pixels <= 8'b01101100;
		12'd3437: row_of_pixels <= 8'b01101100;
		12'd3438: row_of_pixels <= 8'b01101100;
		12'd3439: row_of_pixels <= 8'b01101100;
		12'd3440: row_of_pixels <= 8'b01101100;
		12'd3441: row_of_pixels <= 8'b01101100;
		12'd3442: row_of_pixels <= 8'b01101100;
		12'd3443: row_of_pixels <= 8'b01101100;
		12'd3444: row_of_pixels <= 8'b01101100;
		12'd3445: row_of_pixels <= 8'b01101100;
		12'd3446: row_of_pixels <= 8'b01101100;
		12'd3447: row_of_pixels <= 8'b11111111;
		12'd3448: row_of_pixels <= 8'b01101100;
		12'd3449: row_of_pixels <= 8'b01101100;
		12'd3450: row_of_pixels <= 8'b01101100;
		12'd3451: row_of_pixels <= 8'b01101100;
		12'd3452: row_of_pixels <= 8'b01101100;
		12'd3453: row_of_pixels <= 8'b01101100;
		12'd3454: row_of_pixels <= 8'b01101100;
		12'd3455: row_of_pixels <= 8'b01101100;
		12'd3456: row_of_pixels <= 8'b00011000;
		12'd3457: row_of_pixels <= 8'b00011000;
		12'd3458: row_of_pixels <= 8'b00011000;
		12'd3459: row_of_pixels <= 8'b00011000;
		12'd3460: row_of_pixels <= 8'b00011000;
		12'd3461: row_of_pixels <= 8'b11111111;
		12'd3462: row_of_pixels <= 8'b00011000;
		12'd3463: row_of_pixels <= 8'b11111111;
		12'd3464: row_of_pixels <= 8'b00011000;
		12'd3465: row_of_pixels <= 8'b00011000;
		12'd3466: row_of_pixels <= 8'b00011000;
		12'd3467: row_of_pixels <= 8'b00011000;
		12'd3468: row_of_pixels <= 8'b00011000;
		12'd3469: row_of_pixels <= 8'b00011000;
		12'd3470: row_of_pixels <= 8'b00011000;
		12'd3471: row_of_pixels <= 8'b00011000;
		12'd3472: row_of_pixels <= 8'b00011000;
		12'd3473: row_of_pixels <= 8'b00011000;
		12'd3474: row_of_pixels <= 8'b00011000;
		12'd3475: row_of_pixels <= 8'b00011000;
		12'd3476: row_of_pixels <= 8'b00011000;
		12'd3477: row_of_pixels <= 8'b00011000;
		12'd3478: row_of_pixels <= 8'b00011000;
		12'd3479: row_of_pixels <= 8'b00011111;
		12'd3480: row_of_pixels <= 8'b00000000;
		12'd3481: row_of_pixels <= 8'b00000000;
		12'd3482: row_of_pixels <= 8'b00000000;
		12'd3483: row_of_pixels <= 8'b00000000;
		12'd3484: row_of_pixels <= 8'b00000000;
		12'd3485: row_of_pixels <= 8'b00000000;
		12'd3486: row_of_pixels <= 8'b00000000;
		12'd3487: row_of_pixels <= 8'b00000000;
		12'd3488: row_of_pixels <= 8'b00000000;
		12'd3489: row_of_pixels <= 8'b00000000;
		12'd3490: row_of_pixels <= 8'b00000000;
		12'd3491: row_of_pixels <= 8'b00000000;
		12'd3492: row_of_pixels <= 8'b00000000;
		12'd3493: row_of_pixels <= 8'b00000000;
		12'd3494: row_of_pixels <= 8'b00000000;
		12'd3495: row_of_pixels <= 8'b11111000;
		12'd3496: row_of_pixels <= 8'b00011000;
		12'd3497: row_of_pixels <= 8'b00011000;
		12'd3498: row_of_pixels <= 8'b00011000;
		12'd3499: row_of_pixels <= 8'b00011000;
		12'd3500: row_of_pixels <= 8'b00011000;
		12'd3501: row_of_pixels <= 8'b00011000;
		12'd3502: row_of_pixels <= 8'b00011000;
		12'd3503: row_of_pixels <= 8'b00011000;
		12'd3504: row_of_pixels <= 8'b11111111;
		12'd3505: row_of_pixels <= 8'b11111111;
		12'd3506: row_of_pixels <= 8'b11111111;
		12'd3507: row_of_pixels <= 8'b11111111;
		12'd3508: row_of_pixels <= 8'b11111111;
		12'd3509: row_of_pixels <= 8'b11111111;
		12'd3510: row_of_pixels <= 8'b11111111;
		12'd3511: row_of_pixels <= 8'b11111111;
		12'd3512: row_of_pixels <= 8'b11111111;
		12'd3513: row_of_pixels <= 8'b11111111;
		12'd3514: row_of_pixels <= 8'b11111111;
		12'd3515: row_of_pixels <= 8'b11111111;
		12'd3516: row_of_pixels <= 8'b11111111;
		12'd3517: row_of_pixels <= 8'b11111111;
		12'd3518: row_of_pixels <= 8'b11111111;
		12'd3519: row_of_pixels <= 8'b11111111;
		12'd3520: row_of_pixels <= 8'b00000000;
		12'd3521: row_of_pixels <= 8'b00000000;
		12'd3522: row_of_pixels <= 8'b00000000;
		12'd3523: row_of_pixels <= 8'b00000000;
		12'd3524: row_of_pixels <= 8'b00000000;
		12'd3525: row_of_pixels <= 8'b00000000;
		12'd3526: row_of_pixels <= 8'b00000000;
		12'd3527: row_of_pixels <= 8'b11111111;
		12'd3528: row_of_pixels <= 8'b11111111;
		12'd3529: row_of_pixels <= 8'b11111111;
		12'd3530: row_of_pixels <= 8'b11111111;
		12'd3531: row_of_pixels <= 8'b11111111;
		12'd3532: row_of_pixels <= 8'b11111111;
		12'd3533: row_of_pixels <= 8'b11111111;
		12'd3534: row_of_pixels <= 8'b11111111;
		12'd3535: row_of_pixels <= 8'b11111111;
		12'd3536: row_of_pixels <= 8'b00001111;
		12'd3537: row_of_pixels <= 8'b00001111;
		12'd3538: row_of_pixels <= 8'b00001111;
		12'd3539: row_of_pixels <= 8'b00001111;
		12'd3540: row_of_pixels <= 8'b00001111;
		12'd3541: row_of_pixels <= 8'b00001111;
		12'd3542: row_of_pixels <= 8'b00001111;
		12'd3543: row_of_pixels <= 8'b00001111;
		12'd3544: row_of_pixels <= 8'b00001111;
		12'd3545: row_of_pixels <= 8'b00001111;
		12'd3546: row_of_pixels <= 8'b00001111;
		12'd3547: row_of_pixels <= 8'b00001111;
		12'd3548: row_of_pixels <= 8'b00001111;
		12'd3549: row_of_pixels <= 8'b00001111;
		12'd3550: row_of_pixels <= 8'b00001111;
		12'd3551: row_of_pixels <= 8'b00001111;
		12'd3552: row_of_pixels <= 8'b11110000;
		12'd3553: row_of_pixels <= 8'b11110000;
		12'd3554: row_of_pixels <= 8'b11110000;
		12'd3555: row_of_pixels <= 8'b11110000;
		12'd3556: row_of_pixels <= 8'b11110000;
		12'd3557: row_of_pixels <= 8'b11110000;
		12'd3558: row_of_pixels <= 8'b11110000;
		12'd3559: row_of_pixels <= 8'b11110000;
		12'd3560: row_of_pixels <= 8'b11110000;
		12'd3561: row_of_pixels <= 8'b11110000;
		12'd3562: row_of_pixels <= 8'b11110000;
		12'd3563: row_of_pixels <= 8'b11110000;
		12'd3564: row_of_pixels <= 8'b11110000;
		12'd3565: row_of_pixels <= 8'b11110000;
		12'd3566: row_of_pixels <= 8'b11110000;
		12'd3567: row_of_pixels <= 8'b11110000;
		12'd3568: row_of_pixels <= 8'b11111111;
		12'd3569: row_of_pixels <= 8'b11111111;
		12'd3570: row_of_pixels <= 8'b11111111;
		12'd3571: row_of_pixels <= 8'b11111111;
		12'd3572: row_of_pixels <= 8'b11111111;
		12'd3573: row_of_pixels <= 8'b11111111;
		12'd3574: row_of_pixels <= 8'b11111111;
		12'd3575: row_of_pixels <= 8'b00000000;
		12'd3576: row_of_pixels <= 8'b00000000;
		12'd3577: row_of_pixels <= 8'b00000000;
		12'd3578: row_of_pixels <= 8'b00000000;
		12'd3579: row_of_pixels <= 8'b00000000;
		12'd3580: row_of_pixels <= 8'b00000000;
		12'd3581: row_of_pixels <= 8'b00000000;
		12'd3582: row_of_pixels <= 8'b00000000;
		12'd3583: row_of_pixels <= 8'b00000000;
		12'd3584: row_of_pixels <= 8'b00000000;
		12'd3585: row_of_pixels <= 8'b00000000;
		12'd3586: row_of_pixels <= 8'b00000000;
		12'd3587: row_of_pixels <= 8'b00000000;
		12'd3588: row_of_pixels <= 8'b00000000;
		12'd3589: row_of_pixels <= 8'b01101110;
		12'd3590: row_of_pixels <= 8'b00111011;
		12'd3591: row_of_pixels <= 8'b00011011;
		12'd3592: row_of_pixels <= 8'b00011011;
		12'd3593: row_of_pixels <= 8'b00011011;
		12'd3594: row_of_pixels <= 8'b00111011;
		12'd3595: row_of_pixels <= 8'b01101110;
		12'd3596: row_of_pixels <= 8'b00000000;
		12'd3597: row_of_pixels <= 8'b00000000;
		12'd3598: row_of_pixels <= 8'b00000000;
		12'd3599: row_of_pixels <= 8'b00000000;
		12'd3600: row_of_pixels <= 8'b00000000;
		12'd3601: row_of_pixels <= 8'b00000000;
		12'd3602: row_of_pixels <= 8'b00011110;
		12'd3603: row_of_pixels <= 8'b00110011;
		12'd3604: row_of_pixels <= 8'b00110011;
		12'd3605: row_of_pixels <= 8'b00110011;
		12'd3606: row_of_pixels <= 8'b00011011;
		12'd3607: row_of_pixels <= 8'b00110011;
		12'd3608: row_of_pixels <= 8'b01100011;
		12'd3609: row_of_pixels <= 8'b01100011;
		12'd3610: row_of_pixels <= 8'b01100011;
		12'd3611: row_of_pixels <= 8'b00110011;
		12'd3612: row_of_pixels <= 8'b00000000;
		12'd3613: row_of_pixels <= 8'b00000000;
		12'd3614: row_of_pixels <= 8'b00000000;
		12'd3615: row_of_pixels <= 8'b00000000;
		12'd3616: row_of_pixels <= 8'b00000000;
		12'd3617: row_of_pixels <= 8'b00000000;
		12'd3618: row_of_pixels <= 8'b01111111;
		12'd3619: row_of_pixels <= 8'b01100011;
		12'd3620: row_of_pixels <= 8'b01100011;
		12'd3621: row_of_pixels <= 8'b00000011;
		12'd3622: row_of_pixels <= 8'b00000011;
		12'd3623: row_of_pixels <= 8'b00000011;
		12'd3624: row_of_pixels <= 8'b00000011;
		12'd3625: row_of_pixels <= 8'b00000011;
		12'd3626: row_of_pixels <= 8'b00000011;
		12'd3627: row_of_pixels <= 8'b00000011;
		12'd3628: row_of_pixels <= 8'b00000000;
		12'd3629: row_of_pixels <= 8'b00000000;
		12'd3630: row_of_pixels <= 8'b00000000;
		12'd3631: row_of_pixels <= 8'b00000000;
		12'd3632: row_of_pixels <= 8'b00000000;
		12'd3633: row_of_pixels <= 8'b00000000;
		12'd3634: row_of_pixels <= 8'b00000000;
		12'd3635: row_of_pixels <= 8'b00000000;
		12'd3636: row_of_pixels <= 8'b01111111;
		12'd3637: row_of_pixels <= 8'b00110110;
		12'd3638: row_of_pixels <= 8'b00110110;
		12'd3639: row_of_pixels <= 8'b00110110;
		12'd3640: row_of_pixels <= 8'b00110110;
		12'd3641: row_of_pixels <= 8'b00110110;
		12'd3642: row_of_pixels <= 8'b00110110;
		12'd3643: row_of_pixels <= 8'b00110110;
		12'd3644: row_of_pixels <= 8'b00000000;
		12'd3645: row_of_pixels <= 8'b00000000;
		12'd3646: row_of_pixels <= 8'b00000000;
		12'd3647: row_of_pixels <= 8'b00000000;
		12'd3648: row_of_pixels <= 8'b00000000;
		12'd3649: row_of_pixels <= 8'b00000000;
		12'd3650: row_of_pixels <= 8'b00000000;
		12'd3651: row_of_pixels <= 8'b01111111;
		12'd3652: row_of_pixels <= 8'b01100011;
		12'd3653: row_of_pixels <= 8'b00000110;
		12'd3654: row_of_pixels <= 8'b00001100;
		12'd3655: row_of_pixels <= 8'b00011000;
		12'd3656: row_of_pixels <= 8'b00001100;
		12'd3657: row_of_pixels <= 8'b00000110;
		12'd3658: row_of_pixels <= 8'b01100011;
		12'd3659: row_of_pixels <= 8'b01111111;
		12'd3660: row_of_pixels <= 8'b00000000;
		12'd3661: row_of_pixels <= 8'b00000000;
		12'd3662: row_of_pixels <= 8'b00000000;
		12'd3663: row_of_pixels <= 8'b00000000;
		12'd3664: row_of_pixels <= 8'b00000000;
		12'd3665: row_of_pixels <= 8'b00000000;
		12'd3666: row_of_pixels <= 8'b00000000;
		12'd3667: row_of_pixels <= 8'b00000000;
		12'd3668: row_of_pixels <= 8'b00000000;
		12'd3669: row_of_pixels <= 8'b01111110;
		12'd3670: row_of_pixels <= 8'b00011011;
		12'd3671: row_of_pixels <= 8'b00011011;
		12'd3672: row_of_pixels <= 8'b00011011;
		12'd3673: row_of_pixels <= 8'b00011011;
		12'd3674: row_of_pixels <= 8'b00011011;
		12'd3675: row_of_pixels <= 8'b00001110;
		12'd3676: row_of_pixels <= 8'b00000000;
		12'd3677: row_of_pixels <= 8'b00000000;
		12'd3678: row_of_pixels <= 8'b00000000;
		12'd3679: row_of_pixels <= 8'b00000000;
		12'd3680: row_of_pixels <= 8'b00000000;
		12'd3681: row_of_pixels <= 8'b00000000;
		12'd3682: row_of_pixels <= 8'b00000000;
		12'd3683: row_of_pixels <= 8'b00000000;
		12'd3684: row_of_pixels <= 8'b01100110;
		12'd3685: row_of_pixels <= 8'b01100110;
		12'd3686: row_of_pixels <= 8'b01100110;
		12'd3687: row_of_pixels <= 8'b01100110;
		12'd3688: row_of_pixels <= 8'b01100110;
		12'd3689: row_of_pixels <= 8'b00111110;
		12'd3690: row_of_pixels <= 8'b00000110;
		12'd3691: row_of_pixels <= 8'b00000110;
		12'd3692: row_of_pixels <= 8'b00000011;
		12'd3693: row_of_pixels <= 8'b00000000;
		12'd3694: row_of_pixels <= 8'b00000000;
		12'd3695: row_of_pixels <= 8'b00000000;
		12'd3696: row_of_pixels <= 8'b00000000;
		12'd3697: row_of_pixels <= 8'b00000000;
		12'd3698: row_of_pixels <= 8'b00000000;
		12'd3699: row_of_pixels <= 8'b00000000;
		12'd3700: row_of_pixels <= 8'b01101110;
		12'd3701: row_of_pixels <= 8'b00111011;
		12'd3702: row_of_pixels <= 8'b00011000;
		12'd3703: row_of_pixels <= 8'b00011000;
		12'd3704: row_of_pixels <= 8'b00011000;
		12'd3705: row_of_pixels <= 8'b00011000;
		12'd3706: row_of_pixels <= 8'b00011000;
		12'd3707: row_of_pixels <= 8'b00011000;
		12'd3708: row_of_pixels <= 8'b00000000;
		12'd3709: row_of_pixels <= 8'b00000000;
		12'd3710: row_of_pixels <= 8'b00000000;
		12'd3711: row_of_pixels <= 8'b00000000;
		12'd3712: row_of_pixels <= 8'b00000000;
		12'd3713: row_of_pixels <= 8'b00000000;
		12'd3714: row_of_pixels <= 8'b00000000;
		12'd3715: row_of_pixels <= 8'b01111110;
		12'd3716: row_of_pixels <= 8'b00011000;
		12'd3717: row_of_pixels <= 8'b00111100;
		12'd3718: row_of_pixels <= 8'b01100110;
		12'd3719: row_of_pixels <= 8'b01100110;
		12'd3720: row_of_pixels <= 8'b01100110;
		12'd3721: row_of_pixels <= 8'b00111100;
		12'd3722: row_of_pixels <= 8'b00011000;
		12'd3723: row_of_pixels <= 8'b01111110;
		12'd3724: row_of_pixels <= 8'b00000000;
		12'd3725: row_of_pixels <= 8'b00000000;
		12'd3726: row_of_pixels <= 8'b00000000;
		12'd3727: row_of_pixels <= 8'b00000000;
		12'd3728: row_of_pixels <= 8'b00000000;
		12'd3729: row_of_pixels <= 8'b00000000;
		12'd3730: row_of_pixels <= 8'b00000000;
		12'd3731: row_of_pixels <= 8'b00011100;
		12'd3732: row_of_pixels <= 8'b00110110;
		12'd3733: row_of_pixels <= 8'b01100011;
		12'd3734: row_of_pixels <= 8'b01100011;
		12'd3735: row_of_pixels <= 8'b01111111;
		12'd3736: row_of_pixels <= 8'b01100011;
		12'd3737: row_of_pixels <= 8'b01100011;
		12'd3738: row_of_pixels <= 8'b00110110;
		12'd3739: row_of_pixels <= 8'b00011100;
		12'd3740: row_of_pixels <= 8'b00000000;
		12'd3741: row_of_pixels <= 8'b00000000;
		12'd3742: row_of_pixels <= 8'b00000000;
		12'd3743: row_of_pixels <= 8'b00000000;
		12'd3744: row_of_pixels <= 8'b00000000;
		12'd3745: row_of_pixels <= 8'b00000000;
		12'd3746: row_of_pixels <= 8'b00011100;
		12'd3747: row_of_pixels <= 8'b00110110;
		12'd3748: row_of_pixels <= 8'b01100011;
		12'd3749: row_of_pixels <= 8'b01100011;
		12'd3750: row_of_pixels <= 8'b01100011;
		12'd3751: row_of_pixels <= 8'b00110110;
		12'd3752: row_of_pixels <= 8'b00110110;
		12'd3753: row_of_pixels <= 8'b00110110;
		12'd3754: row_of_pixels <= 8'b00110110;
		12'd3755: row_of_pixels <= 8'b01110111;
		12'd3756: row_of_pixels <= 8'b00000000;
		12'd3757: row_of_pixels <= 8'b00000000;
		12'd3758: row_of_pixels <= 8'b00000000;
		12'd3759: row_of_pixels <= 8'b00000000;
		12'd3760: row_of_pixels <= 8'b00000000;
		12'd3761: row_of_pixels <= 8'b00000000;
		12'd3762: row_of_pixels <= 8'b01111000;
		12'd3763: row_of_pixels <= 8'b00001100;
		12'd3764: row_of_pixels <= 8'b00011000;
		12'd3765: row_of_pixels <= 8'b00110000;
		12'd3766: row_of_pixels <= 8'b01111100;
		12'd3767: row_of_pixels <= 8'b01100110;
		12'd3768: row_of_pixels <= 8'b01100110;
		12'd3769: row_of_pixels <= 8'b01100110;
		12'd3770: row_of_pixels <= 8'b01100110;
		12'd3771: row_of_pixels <= 8'b00111100;
		12'd3772: row_of_pixels <= 8'b00000000;
		12'd3773: row_of_pixels <= 8'b00000000;
		12'd3774: row_of_pixels <= 8'b00000000;
		12'd3775: row_of_pixels <= 8'b00000000;
		12'd3776: row_of_pixels <= 8'b00000000;
		12'd3777: row_of_pixels <= 8'b00000000;
		12'd3778: row_of_pixels <= 8'b00000000;
		12'd3779: row_of_pixels <= 8'b00000000;
		12'd3780: row_of_pixels <= 8'b00000000;
		12'd3781: row_of_pixels <= 8'b01111110;
		12'd3782: row_of_pixels <= 8'b11011011;
		12'd3783: row_of_pixels <= 8'b11011011;
		12'd3784: row_of_pixels <= 8'b11011011;
		12'd3785: row_of_pixels <= 8'b01111110;
		12'd3786: row_of_pixels <= 8'b00000000;
		12'd3787: row_of_pixels <= 8'b00000000;
		12'd3788: row_of_pixels <= 8'b00000000;
		12'd3789: row_of_pixels <= 8'b00000000;
		12'd3790: row_of_pixels <= 8'b00000000;
		12'd3791: row_of_pixels <= 8'b00000000;
		12'd3792: row_of_pixels <= 8'b00000000;
		12'd3793: row_of_pixels <= 8'b00000000;
		12'd3794: row_of_pixels <= 8'b00000000;
		12'd3795: row_of_pixels <= 8'b11000000;
		12'd3796: row_of_pixels <= 8'b01100000;
		12'd3797: row_of_pixels <= 8'b01111110;
		12'd3798: row_of_pixels <= 8'b11011011;
		12'd3799: row_of_pixels <= 8'b11011011;
		12'd3800: row_of_pixels <= 8'b11001111;
		12'd3801: row_of_pixels <= 8'b01111110;
		12'd3802: row_of_pixels <= 8'b00000110;
		12'd3803: row_of_pixels <= 8'b00000011;
		12'd3804: row_of_pixels <= 8'b00000000;
		12'd3805: row_of_pixels <= 8'b00000000;
		12'd3806: row_of_pixels <= 8'b00000000;
		12'd3807: row_of_pixels <= 8'b00000000;
		12'd3808: row_of_pixels <= 8'b00000000;
		12'd3809: row_of_pixels <= 8'b00000000;
		12'd3810: row_of_pixels <= 8'b00111000;
		12'd3811: row_of_pixels <= 8'b00001100;
		12'd3812: row_of_pixels <= 8'b00000110;
		12'd3813: row_of_pixels <= 8'b00000110;
		12'd3814: row_of_pixels <= 8'b00111110;
		12'd3815: row_of_pixels <= 8'b00000110;
		12'd3816: row_of_pixels <= 8'b00000110;
		12'd3817: row_of_pixels <= 8'b00000110;
		12'd3818: row_of_pixels <= 8'b00001100;
		12'd3819: row_of_pixels <= 8'b00111000;
		12'd3820: row_of_pixels <= 8'b00000000;
		12'd3821: row_of_pixels <= 8'b00000000;
		12'd3822: row_of_pixels <= 8'b00000000;
		12'd3823: row_of_pixels <= 8'b00000000;
		12'd3824: row_of_pixels <= 8'b00000000;
		12'd3825: row_of_pixels <= 8'b00000000;
		12'd3826: row_of_pixels <= 8'b00000000;
		12'd3827: row_of_pixels <= 8'b00111110;
		12'd3828: row_of_pixels <= 8'b01100011;
		12'd3829: row_of_pixels <= 8'b01100011;
		12'd3830: row_of_pixels <= 8'b01100011;
		12'd3831: row_of_pixels <= 8'b01100011;
		12'd3832: row_of_pixels <= 8'b01100011;
		12'd3833: row_of_pixels <= 8'b01100011;
		12'd3834: row_of_pixels <= 8'b01100011;
		12'd3835: row_of_pixels <= 8'b01100011;
		12'd3836: row_of_pixels <= 8'b00000000;
		12'd3837: row_of_pixels <= 8'b00000000;
		12'd3838: row_of_pixels <= 8'b00000000;
		12'd3839: row_of_pixels <= 8'b00000000;
		12'd3840: row_of_pixels <= 8'b00000000;
		12'd3841: row_of_pixels <= 8'b00000000;
		12'd3842: row_of_pixels <= 8'b00000000;
		12'd3843: row_of_pixels <= 8'b00000000;
		12'd3844: row_of_pixels <= 8'b01111111;
		12'd3845: row_of_pixels <= 8'b00000000;
		12'd3846: row_of_pixels <= 8'b00000000;
		12'd3847: row_of_pixels <= 8'b01111111;
		12'd3848: row_of_pixels <= 8'b00000000;
		12'd3849: row_of_pixels <= 8'b00000000;
		12'd3850: row_of_pixels <= 8'b01111111;
		12'd3851: row_of_pixels <= 8'b00000000;
		12'd3852: row_of_pixels <= 8'b00000000;
		12'd3853: row_of_pixels <= 8'b00000000;
		12'd3854: row_of_pixels <= 8'b00000000;
		12'd3855: row_of_pixels <= 8'b00000000;
		12'd3856: row_of_pixels <= 8'b00000000;
		12'd3857: row_of_pixels <= 8'b00000000;
		12'd3858: row_of_pixels <= 8'b00000000;
		12'd3859: row_of_pixels <= 8'b00000000;
		12'd3860: row_of_pixels <= 8'b00011000;
		12'd3861: row_of_pixels <= 8'b00011000;
		12'd3862: row_of_pixels <= 8'b01111110;
		12'd3863: row_of_pixels <= 8'b00011000;
		12'd3864: row_of_pixels <= 8'b00011000;
		12'd3865: row_of_pixels <= 8'b00000000;
		12'd3866: row_of_pixels <= 8'b00000000;
		12'd3867: row_of_pixels <= 8'b11111111;
		12'd3868: row_of_pixels <= 8'b00000000;
		12'd3869: row_of_pixels <= 8'b00000000;
		12'd3870: row_of_pixels <= 8'b00000000;
		12'd3871: row_of_pixels <= 8'b00000000;
		12'd3872: row_of_pixels <= 8'b00000000;
		12'd3873: row_of_pixels <= 8'b00000000;
		12'd3874: row_of_pixels <= 8'b00000000;
		12'd3875: row_of_pixels <= 8'b00001100;
		12'd3876: row_of_pixels <= 8'b00011000;
		12'd3877: row_of_pixels <= 8'b00110000;
		12'd3878: row_of_pixels <= 8'b01100000;
		12'd3879: row_of_pixels <= 8'b00110000;
		12'd3880: row_of_pixels <= 8'b00011000;
		12'd3881: row_of_pixels <= 8'b00001100;
		12'd3882: row_of_pixels <= 8'b00000000;
		12'd3883: row_of_pixels <= 8'b01111110;
		12'd3884: row_of_pixels <= 8'b00000000;
		12'd3885: row_of_pixels <= 8'b00000000;
		12'd3886: row_of_pixels <= 8'b00000000;
		12'd3887: row_of_pixels <= 8'b00000000;
		12'd3888: row_of_pixels <= 8'b00000000;
		12'd3889: row_of_pixels <= 8'b00000000;
		12'd3890: row_of_pixels <= 8'b00000000;
		12'd3891: row_of_pixels <= 8'b00110000;
		12'd3892: row_of_pixels <= 8'b00011000;
		12'd3893: row_of_pixels <= 8'b00001100;
		12'd3894: row_of_pixels <= 8'b00000110;
		12'd3895: row_of_pixels <= 8'b00001100;
		12'd3896: row_of_pixels <= 8'b00011000;
		12'd3897: row_of_pixels <= 8'b00110000;
		12'd3898: row_of_pixels <= 8'b00000000;
		12'd3899: row_of_pixels <= 8'b01111110;
		12'd3900: row_of_pixels <= 8'b00000000;
		12'd3901: row_of_pixels <= 8'b00000000;
		12'd3902: row_of_pixels <= 8'b00000000;
		12'd3903: row_of_pixels <= 8'b00000000;
		12'd3904: row_of_pixels <= 8'b00000000;
		12'd3905: row_of_pixels <= 8'b00000000;
		12'd3906: row_of_pixels <= 8'b01110000;
		12'd3907: row_of_pixels <= 8'b11011000;
		12'd3908: row_of_pixels <= 8'b11011000;
		12'd3909: row_of_pixels <= 8'b11011000;
		12'd3910: row_of_pixels <= 8'b00011000;
		12'd3911: row_of_pixels <= 8'b00011000;
		12'd3912: row_of_pixels <= 8'b00011000;
		12'd3913: row_of_pixels <= 8'b00011000;
		12'd3914: row_of_pixels <= 8'b00011000;
		12'd3915: row_of_pixels <= 8'b00011000;
		12'd3916: row_of_pixels <= 8'b00011000;
		12'd3917: row_of_pixels <= 8'b00011000;
		12'd3918: row_of_pixels <= 8'b00011000;
		12'd3919: row_of_pixels <= 8'b00011000;
		12'd3920: row_of_pixels <= 8'b00011000;
		12'd3921: row_of_pixels <= 8'b00011000;
		12'd3922: row_of_pixels <= 8'b00011000;
		12'd3923: row_of_pixels <= 8'b00011000;
		12'd3924: row_of_pixels <= 8'b00011000;
		12'd3925: row_of_pixels <= 8'b00011000;
		12'd3926: row_of_pixels <= 8'b00011000;
		12'd3927: row_of_pixels <= 8'b00011000;
		12'd3928: row_of_pixels <= 8'b00011011;
		12'd3929: row_of_pixels <= 8'b00011011;
		12'd3930: row_of_pixels <= 8'b00011011;
		12'd3931: row_of_pixels <= 8'b00001110;
		12'd3932: row_of_pixels <= 8'b00000000;
		12'd3933: row_of_pixels <= 8'b00000000;
		12'd3934: row_of_pixels <= 8'b00000000;
		12'd3935: row_of_pixels <= 8'b00000000;
		12'd3936: row_of_pixels <= 8'b00000000;
		12'd3937: row_of_pixels <= 8'b00000000;
		12'd3938: row_of_pixels <= 8'b00000000;
		12'd3939: row_of_pixels <= 8'b00000000;
		12'd3940: row_of_pixels <= 8'b00011000;
		12'd3941: row_of_pixels <= 8'b00011000;
		12'd3942: row_of_pixels <= 8'b00000000;
		12'd3943: row_of_pixels <= 8'b01111110;
		12'd3944: row_of_pixels <= 8'b00000000;
		12'd3945: row_of_pixels <= 8'b00011000;
		12'd3946: row_of_pixels <= 8'b00011000;
		12'd3947: row_of_pixels <= 8'b00000000;
		12'd3948: row_of_pixels <= 8'b00000000;
		12'd3949: row_of_pixels <= 8'b00000000;
		12'd3950: row_of_pixels <= 8'b00000000;
		12'd3951: row_of_pixels <= 8'b00000000;
		12'd3952: row_of_pixels <= 8'b00000000;
		12'd3953: row_of_pixels <= 8'b00000000;
		12'd3954: row_of_pixels <= 8'b00000000;
		12'd3955: row_of_pixels <= 8'b00000000;
		12'd3956: row_of_pixels <= 8'b00000000;
		12'd3957: row_of_pixels <= 8'b01101110;
		12'd3958: row_of_pixels <= 8'b00111011;
		12'd3959: row_of_pixels <= 8'b00000000;
		12'd3960: row_of_pixels <= 8'b01101110;
		12'd3961: row_of_pixels <= 8'b00111011;
		12'd3962: row_of_pixels <= 8'b00000000;
		12'd3963: row_of_pixels <= 8'b00000000;
		12'd3964: row_of_pixels <= 8'b00000000;
		12'd3965: row_of_pixels <= 8'b00000000;
		12'd3966: row_of_pixels <= 8'b00000000;
		12'd3967: row_of_pixels <= 8'b00000000;
		12'd3968: row_of_pixels <= 8'b00000000;
		12'd3969: row_of_pixels <= 8'b00011100;
		12'd3970: row_of_pixels <= 8'b00110110;
		12'd3971: row_of_pixels <= 8'b00110110;
		12'd3972: row_of_pixels <= 8'b00011100;
		12'd3973: row_of_pixels <= 8'b00000000;
		12'd3974: row_of_pixels <= 8'b00000000;
		12'd3975: row_of_pixels <= 8'b00000000;
		12'd3976: row_of_pixels <= 8'b00000000;
		12'd3977: row_of_pixels <= 8'b00000000;
		12'd3978: row_of_pixels <= 8'b00000000;
		12'd3979: row_of_pixels <= 8'b00000000;
		12'd3980: row_of_pixels <= 8'b00000000;
		12'd3981: row_of_pixels <= 8'b00000000;
		12'd3982: row_of_pixels <= 8'b00000000;
		12'd3983: row_of_pixels <= 8'b00000000;
		12'd3984: row_of_pixels <= 8'b00000000;
		12'd3985: row_of_pixels <= 8'b00000000;
		12'd3986: row_of_pixels <= 8'b00000000;
		12'd3987: row_of_pixels <= 8'b00000000;
		12'd3988: row_of_pixels <= 8'b00000000;
		12'd3989: row_of_pixels <= 8'b00000000;
		12'd3990: row_of_pixels <= 8'b00000000;
		12'd3991: row_of_pixels <= 8'b00011000;
		12'd3992: row_of_pixels <= 8'b00011000;
		12'd3993: row_of_pixels <= 8'b00000000;
		12'd3994: row_of_pixels <= 8'b00000000;
		12'd3995: row_of_pixels <= 8'b00000000;
		12'd3996: row_of_pixels <= 8'b00000000;
		12'd3997: row_of_pixels <= 8'b00000000;
		12'd3998: row_of_pixels <= 8'b00000000;
		12'd3999: row_of_pixels <= 8'b00000000;
		12'd4000: row_of_pixels <= 8'b00000000;
		12'd4001: row_of_pixels <= 8'b00000000;
		12'd4002: row_of_pixels <= 8'b00000000;
		12'd4003: row_of_pixels <= 8'b00000000;
		12'd4004: row_of_pixels <= 8'b00000000;
		12'd4005: row_of_pixels <= 8'b00000000;
		12'd4006: row_of_pixels <= 8'b00000000;
		12'd4007: row_of_pixels <= 8'b00000000;
		12'd4008: row_of_pixels <= 8'b00011000;
		12'd4009: row_of_pixels <= 8'b00000000;
		12'd4010: row_of_pixels <= 8'b00000000;
		12'd4011: row_of_pixels <= 8'b00000000;
		12'd4012: row_of_pixels <= 8'b00000000;
		12'd4013: row_of_pixels <= 8'b00000000;
		12'd4014: row_of_pixels <= 8'b00000000;
		12'd4015: row_of_pixels <= 8'b00000000;
		12'd4016: row_of_pixels <= 8'b00000000;
		12'd4017: row_of_pixels <= 8'b11110000;
		12'd4018: row_of_pixels <= 8'b00110000;
		12'd4019: row_of_pixels <= 8'b00110000;
		12'd4020: row_of_pixels <= 8'b00110000;
		12'd4021: row_of_pixels <= 8'b00110000;
		12'd4022: row_of_pixels <= 8'b00110000;
		12'd4023: row_of_pixels <= 8'b00110111;
		12'd4024: row_of_pixels <= 8'b00110110;
		12'd4025: row_of_pixels <= 8'b00110110;
		12'd4026: row_of_pixels <= 8'b00111100;
		12'd4027: row_of_pixels <= 8'b00111000;
		12'd4028: row_of_pixels <= 8'b00000000;
		12'd4029: row_of_pixels <= 8'b00000000;
		12'd4030: row_of_pixels <= 8'b00000000;
		12'd4031: row_of_pixels <= 8'b00000000;
		12'd4032: row_of_pixels <= 8'b00000000;
		12'd4033: row_of_pixels <= 8'b00011011;
		12'd4034: row_of_pixels <= 8'b00110110;
		12'd4035: row_of_pixels <= 8'b00110110;
		12'd4036: row_of_pixels <= 8'b00110110;
		12'd4037: row_of_pixels <= 8'b00110110;
		12'd4038: row_of_pixels <= 8'b00110110;
		12'd4039: row_of_pixels <= 8'b00000000;
		12'd4040: row_of_pixels <= 8'b00000000;
		12'd4041: row_of_pixels <= 8'b00000000;
		12'd4042: row_of_pixels <= 8'b00000000;
		12'd4043: row_of_pixels <= 8'b00000000;
		12'd4044: row_of_pixels <= 8'b00000000;
		12'd4045: row_of_pixels <= 8'b00000000;
		12'd4046: row_of_pixels <= 8'b00000000;
		12'd4047: row_of_pixels <= 8'b00000000;
		12'd4048: row_of_pixels <= 8'b00000000;
		12'd4049: row_of_pixels <= 8'b00001110;
		12'd4050: row_of_pixels <= 8'b00011011;
		12'd4051: row_of_pixels <= 8'b00001100;
		12'd4052: row_of_pixels <= 8'b00000110;
		12'd4053: row_of_pixels <= 8'b00010011;
		12'd4054: row_of_pixels <= 8'b00011111;
		12'd4055: row_of_pixels <= 8'b00000000;
		12'd4056: row_of_pixels <= 8'b00000000;
		12'd4057: row_of_pixels <= 8'b00000000;
		12'd4058: row_of_pixels <= 8'b00000000;
		12'd4059: row_of_pixels <= 8'b00000000;
		12'd4060: row_of_pixels <= 8'b00000000;
		12'd4061: row_of_pixels <= 8'b00000000;
		12'd4062: row_of_pixels <= 8'b00000000;
		12'd4063: row_of_pixels <= 8'b00000000;
		12'd4064: row_of_pixels <= 8'b00000000;
		12'd4065: row_of_pixels <= 8'b00000000;
		12'd4066: row_of_pixels <= 8'b00000000;
		12'd4067: row_of_pixels <= 8'b00000000;
		12'd4068: row_of_pixels <= 8'b00111110;
		12'd4069: row_of_pixels <= 8'b00111110;
		12'd4070: row_of_pixels <= 8'b00111110;
		12'd4071: row_of_pixels <= 8'b00111110;
		12'd4072: row_of_pixels <= 8'b00111110;
		12'd4073: row_of_pixels <= 8'b00111110;
		12'd4074: row_of_pixels <= 8'b00111110;
		12'd4075: row_of_pixels <= 8'b00000000;
		12'd4076: row_of_pixels <= 8'b00000000;
		12'd4077: row_of_pixels <= 8'b00000000;
		12'd4078: row_of_pixels <= 8'b00000000;
		12'd4079: row_of_pixels <= 8'b00000000;
		12'd4080: row_of_pixels <= 8'b00000000;
		12'd4081: row_of_pixels <= 8'b00000000;
		12'd4082: row_of_pixels <= 8'b00000000;
		12'd4083: row_of_pixels <= 8'b00000000;
		12'd4084: row_of_pixels <= 8'b00000000;
		12'd4085: row_of_pixels <= 8'b00000000;
		12'd4086: row_of_pixels <= 8'b00000000;
		12'd4087: row_of_pixels <= 8'b00000000;
		12'd4088: row_of_pixels <= 8'b00000000;
		12'd4089: row_of_pixels <= 8'b00000000;
		12'd4090: row_of_pixels <= 8'b00000000;
		12'd4091: row_of_pixels <= 8'b00000000;
		12'd4092: row_of_pixels <= 8'b00000000;
		12'd4093: row_of_pixels <= 8'b00000000;
		12'd4094: row_of_pixels <= 8'b00000000;
		12'd4095: row_of_pixels <= 8'b00000000;
	endcase
end

endmodule